-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Jul 10 2019 22:39:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    LED1 : out std_logic;
    CLK_3P3_MHZ : in std_logic;
    BTN1 : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__39686\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12023\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_5\ : std_logic;
signal \processor_zipi8.flags_i.un5_shift_carry_value_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.shift_carry_value_1_0_0_cascade_\ : std_logic;
signal \processor_zipi8.stack_i.data_out_ram_0\ : std_logic;
signal \processor_zipi8.shadow_carry_flag\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI88F42_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV3DI8_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIM5NP1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINR4G8_7\ : std_logic;
signal \processor_zipi8.port_id_7_cascade_\ : std_logic;
signal \processor_zipi8.port_id_7\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_7\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_7\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_7_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_7\ : std_logic;
signal \processor_zipi8.stack_memory_5\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_5\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_5_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_5\ : std_logic;
signal \processor_zipi8.port_id_5_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_5\ : std_logic;
signal \processor_zipi8.port_id_5\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_5\ : std_logic;
signal \processor_zipi8.stack_memory_9\ : std_logic;
signal \processor_zipi8.stack_memory_4\ : std_logic;
signal \processor_zipi8.stack_memory_8\ : std_logic;
signal \processor_zipi8.stack_memory_10\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_9\ : std_logic;
signal \processor_zipi8.sy_5\ : std_logic;
signal \processor_zipi8.sy_7\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_8\ : std_logic;
signal \processor_zipi8.pc_vector_8_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_9_cascade_\ : std_logic;
signal address_9 : std_logic;
signal \processor_zipi8.program_counter_i.un380_half_pc_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_10_cascade_\ : std_logic;
signal address_10 : std_logic;
signal \processor_zipi8.return_vector_10\ : std_logic;
signal \processor_zipi8.program_counter_i.un395_half_pcZ0\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_46_7\ : std_logic;
signal \processor_zipi8.pc_vector_8\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_46_7_cascade_\ : std_logic;
signal address_8 : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_8\ : std_logic;
signal \processor_zipi8.flags_i.zero_flag_3_cascade_\ : std_logic;
signal \processor_zipi8.shadow_zero_flag\ : std_logic;
signal \processor_zipi8.alu_result_7\ : std_logic;
signal \processor_zipi8.alu_result_6_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.zero_flag_3_0_5\ : std_logic;
signal \processor_zipi8.alu_result_5\ : std_logic;
signal \processor_zipi8.stack_i.stack_zero_flag\ : std_logic;
signal \processor_zipi8.stack_i.shadow_zero_value\ : std_logic;
signal \processor_zipi8.alu_result_3\ : std_logic;
signal \processor_zipi8.flags_i.m82_1_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.m82_1\ : std_logic;
signal \processor_zipi8.zero_flag_RNIJSPM4\ : std_logic;
signal \processor_zipi8.flags_i.N_55\ : std_logic;
signal \processor_zipi8.flags_i.m61_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIK2TR1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_7\ : std_logic;
signal \processor_zipi8.spm_data_5\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_6\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_6_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_6\ : std_logic;
signal \processor_zipi8.sy_6\ : std_logic;
signal \processor_zipi8.port_id_6_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_6\ : std_logic;
signal \processor_zipi8.port_id_6\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_6\ : std_logic;
signal \processor_zipi8.stack_memory_6\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_6\ : std_logic;
signal \processor_zipi8.flags_i.N_125_mux_cascade_\ : std_logic;
signal \processor_zipi8.stack_i.stack_bit\ : std_logic;
signal \processor_zipi8.run\ : std_logic;
signal \BTN1_c\ : std_logic;
signal \processor_zipi8.stack_memory_2\ : std_logic;
signal \processor_zipi8.special_bit\ : std_logic;
signal \processor_zipi8.state_machine_i.bram_enable\ : std_logic;
signal \processor_zipi8.stack_memory_11\ : std_logic;
signal \processor_zipi8.flags_i.N_37\ : std_logic;
signal \processor_zipi8.stack_memory_7\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_7\ : std_logic;
signal \processor_zipi8.stack_memory_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_155\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_195_cascade_\ : std_logic;
signal address_6 : std_logic;
signal address_4 : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_4\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_4_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_28_4_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_34_5\ : std_logic;
signal \processor_zipi8.pc_vector_6\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_34_5_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_6\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_40_6\ : std_logic;
signal \processor_zipi8.pc_vector_7\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_40_6_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_7\ : std_logic;
signal address_7 : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_5\ : std_logic;
signal \processor_zipi8.pc_vector_5\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_28_4\ : std_logic;
signal address_5 : std_logic;
signal \processor_zipi8.return_vector_11\ : std_logic;
signal \processor_zipi8.program_counter_i.un3_half_pcZ0_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_10\ : std_logic;
signal \processor_zipi8.program_counter_i.un431_half_pc\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_11_cascade_\ : std_logic;
signal \processor_zipi8.address_11\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_9\ : std_logic;
signal \processor_zipi8.pc_vector_9\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_52_8\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_58_9\ : std_logic;
signal \processor_zipi8.flags_i.m49_ns_1\ : std_logic;
signal \processor_zipi8.flags_i.N_50_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.N_51_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.N_123_mux\ : std_logic;
signal \processor_zipi8.flags_i.N_45\ : std_logic;
signal \processor_zipi8.flags_i.m91_amZ0_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.m25_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.N_26_0_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.N_27_0\ : std_logic;
signal \processor_zipi8.flags_i.m20_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.N_21_0\ : std_logic;
signal \processor_zipi8.flags_i.N_1235_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.zero_flag_RNI89VZ0Z91\ : std_logic;
signal \processor_zipi8.flags_i.N_1239\ : std_logic;
signal \processor_zipi8.flags_i.N_124_mux\ : std_logic;
signal \processor_zipi8.flags_i.N_1241_cascade_\ : std_logic;
signal \processor_zipi8.zero_flag_RNIDS654\ : std_logic;
signal \processor_zipi8.stack_pointer_1\ : std_logic;
signal \processor_zipi8.flags_i.m75_amZ0\ : std_logic;
signal \processor_zipi8.flags_i.m75_amZ0_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.zero_flag_RNI3VCZ0Z94\ : std_logic;
signal \processor_zipi8.zero_flag_RNI5GK75\ : std_logic;
signal \processor_zipi8.flags_i.N_1241\ : std_logic;
signal \processor_zipi8.stack_pointer_0\ : std_logic;
signal \processor_zipi8.stack_pointer_2\ : std_logic;
signal \processor_zipi8.flags_i.N_54\ : std_logic;
signal \processor_zipi8.flags_i.m68_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_6\ : std_logic;
signal \processor_zipi8.spm_data_6\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe8\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe11\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212_cascade_\ : std_logic;
signal \processor_zipi8.shift_rotate_result_6\ : std_logic;
signal \processor_zipi8.shift_rotate_result_5\ : std_logic;
signal \processor_zipi8.port_id_2_cascade_\ : std_logic;
signal \processor_zipi8.port_id_2\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_2\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_2\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_2_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_2\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_2\ : std_logic;
signal \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_0_cascade_\ : std_logic;
signal instruction_2 : std_logic;
signal \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_1_cascade_\ : std_logic;
signal \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_0\ : std_logic;
signal address_2 : std_logic;
signal \processor_zipi8.stack_pointer_4\ : std_logic;
signal \processor_zipi8.flags_i.N_34\ : std_logic;
signal \processor_zipi8.port_id_0_cascade_\ : std_logic;
signal \processor_zipi8.stack_memory_0\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_0\ : std_logic;
signal \processor_zipi8.pc_vector_0\ : std_logic;
signal \processor_zipi8.pc_vector_0_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_0\ : std_logic;
signal \processor_zipi8.flags_i.i14_mux\ : std_logic;
signal \processor_zipi8.flags_i.i14_mux_0\ : std_logic;
signal \processor_zipi8.zero_flag_RNIC4FP9\ : std_logic;
signal \processor_zipi8.program_counter_i.t_state_0_1\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_1_cascade_\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_1_cascade_\ : std_logic;
signal address_1 : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0\ : std_logic;
signal address_0 : std_logic;
signal \processor_zipi8.zero_flag_RNIL8RB5\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_1\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_4_0\ : std_logic;
signal \processor_zipi8.program_counter_i.carry_pc_22_3\ : std_logic;
signal \processor_zipi8.pc_vector_2\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_2\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_2\ : std_logic;
signal \processor_zipi8.program_counter_i.un3_half_pcZ0\ : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_3\ : std_logic;
signal \processor_zipi8.un16_alu_mux_sel_value_cascade_\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.un23_flag_enable_type\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_1_cascade_\ : std_logic;
signal \processor_zipi8.shift_rotate_result_2\ : std_logic;
signal \processor_zipi8.spm_data_2\ : std_logic;
signal \processor_zipi8.register_bank_control_i.un31_regbank_type_3_cascade_\ : std_logic;
signal \processor_zipi8.register_bank_control_i.un31_regbank_type\ : std_logic;
signal \processor_zipi8.shift_rotate_result_0\ : std_logic;
signal \processor_zipi8.spm_data_0\ : std_logic;
signal \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_0_cascade_\ : std_logic;
signal \processor_zipi8.pc_mode_2_0_0\ : std_logic;
signal \processor_zipi8.decode4_pc_statck_i.un3_pc_modeZ0\ : std_logic;
signal \processor_zipi8.N_17_0\ : std_logic;
signal bram_enable_g : std_logic;
signal \processor_zipi8.flags_i.m104Z0Z_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI44F42_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIK4HN1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNII1NP1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIGUSR1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7B4G8_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe13\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe15\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe9\ : std_logic;
signal \processor_zipi8.sx_7\ : std_logic;
signal \processor_zipi8.sx_6\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_7\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_6\ : std_logic;
signal \processor_zipi8.flags_i.carry_flag_value_1_1_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.parity_4\ : std_logic;
signal \processor_zipi8.flags_i.carry_flag_RNOZ0Z_1\ : std_logic;
signal \processor_zipi8.flags_i.arith_carryZ0\ : std_logic;
signal \processor_zipi8.flags_i.shift_carryZ0\ : std_logic;
signal \processor_zipi8.flags_i.carry_flag_value_1_0_0\ : std_logic;
signal \processor_zipi8.decode4_pc_statck_i.N_22_0\ : std_logic;
signal \processor_zipi8.register_bank_control_i.un17_regbank_type_1\ : std_logic;
signal \processor_zipi8.flags_i.un17_carry_flag_value_0\ : std_logic;
signal \processor_zipi8.alu_mux_sel_value_1\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_0_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_0_cascade_\ : std_logic;
signal \processor_zipi8.port_id_0\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_0\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4Z0Z_0\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1\ : std_logic;
signal instruction_0 : std_logic;
signal \processor_zipi8.register_bank_control_i.un1_bank_value\ : std_logic;
signal \processor_zipi8.register_bank_control_i.bank_0_1_cascade_\ : std_logic;
signal \processor_zipi8.sy_4\ : std_logic;
signal \processor_zipi8.stack_i.stack_bank\ : std_logic;
signal \processor_zipi8.shadow_bank\ : std_logic;
signal \processor_zipi8.un16_alu_mux_sel_value\ : std_logic;
signal \processor_zipi8.un4_arith_logical_sel_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.carry_flag_value_1_0\ : std_logic;
signal \processor_zipi8.internal_reset\ : std_logic;
signal \processor_zipi8.flags_i.N_69\ : std_logic;
signal \processor_zipi8.stack_pointer_3\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_3_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_3\ : std_logic;
signal \processor_zipi8.port_id_3_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_3\ : std_logic;
signal \processor_zipi8.port_id_3\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_3\ : std_logic;
signal instruction_3 : std_logic;
signal \processor_zipi8.pc_vector_3\ : std_logic;
signal \processor_zipi8.pc_mode_2\ : std_logic;
signal \processor_zipi8.pc_mode_1\ : std_logic;
signal address_3 : std_logic;
signal \processor_zipi8.program_counter_i.half_pc_0_0_3\ : std_logic;
signal \processor_zipi8.arith_carry_in_0\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0\ : std_logic;
signal \processor_zipi8.returni_type_o_2\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_3\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.un9_flag_enable_type_cascade_\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_0_cascade_\ : std_logic;
signal \processor_zipi8.flag_enable\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.spm_enable_value_1\ : std_logic;
signal \processor_zipi8.spm_enable\ : std_logic;
signal \processor_zipi8.flags_i.use_zero_flagZ0\ : std_logic;
signal \processor_zipi8.alu_result_0_cascade_\ : std_logic;
signal \processor_zipi8.zero_flag\ : std_logic;
signal \processor_zipi8.carry_flag\ : std_logic;
signal \processor_zipi8.N_11_0\ : std_logic;
signal \processor_zipi8.alu_result_1\ : std_logic;
signal \processor_zipi8.alu_result_2_cascade_\ : std_logic;
signal \processor_zipi8.flags_i.zero_flag_3_0_0\ : std_logic;
signal \processor_zipi8.flags_i.zero_flag_3_0_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe12\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_bm_1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_179\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_am_1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.shift_rotate_result_4\ : std_logic;
signal \processor_zipi8.spm_data_4\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4\ : std_logic;
signal \processor_zipi8.shift_rotate_result_1\ : std_logic;
signal \processor_zipi8.spm_data_1\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.un8_register_enable_type\ : std_logic;
signal \processor_zipi8.t_state_1\ : std_logic;
signal \processor_zipi8.decode4_strobes_enables_i.register_enable_type_0_cascade_\ : std_logic;
signal instruction_17 : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_22_3\ : std_logic;
signal \processor_zipi8.sx_5\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_34_5\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_5\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4\ : std_logic;
signal \processor_zipi8.flags_i.parity_5\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_1_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tzZ0Z_4\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_4_cascade_\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_4\ : std_logic;
signal \processor_zipi8.port_id_4\ : std_logic;
signal \processor_zipi8.arith_logical_sel_1\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_4\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical\ : std_logic;
signal \processor_zipi8.un4_arith_logical_sel\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1Z0Z_1\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.N_773_tz\ : std_logic;
signal \processor_zipi8.arith_logical_sel_1_0_0\ : std_logic;
signal \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_4\ : std_logic;
signal instruction_14 : std_logic;
signal \processor_zipi8.arith_logical_sel_1_0_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_3\ : std_logic;
signal \processor_zipi8.sy_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_bm_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI8OGN1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_am_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIONE42_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI6LMP1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI4ISR1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINP2G8_3_cascade_\ : std_logic;
signal \processor_zipi8.sx_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6\ : std_logic;
signal \processor_zipi8.alu_result_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI43VU1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIGMK32_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIO8HN1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNICBE42_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIQ8MP1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIO5SR1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI781G8_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209\ : std_logic;
signal \processor_zipi8.register_enable\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNISBGN1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_7\ : std_logic;
signal \processor_zipi8.port_id_1\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_1\ : std_logic;
signal instruction_1 : std_logic;
signal \processor_zipi8.pc_vector_1\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_4\ : std_logic;
signal instruction_12 : std_logic;
signal \processor_zipi8.pc_vector_4\ : std_logic;
signal instruction_13 : std_logic;
signal \processor_zipi8.sx_0\ : std_logic;
signal \LED1_c\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_119_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_95\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_151\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_175\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_191_cascade_\ : std_logic;
signal \processor_zipi8.sx_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNII4IQ1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI4AK32_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIOMUU1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI8MSR1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIAPMP1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFIBI8_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7A3G8_4_cascade_\ : std_logic;
signal \processor_zipi8.sx_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNISRE42_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI4KGN1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIKJE42_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI0ESR1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI2HMP1_2\ : std_logic;
signal \processor_zipi8.sx_addr_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI792G8_2_cascade_\ : std_logic;
signal \processor_zipi8.sx_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_0\ : std_logic;
signal \processor_zipi8.shift_rotate_result_3\ : std_logic;
signal \processor_zipi8.spm_data_3\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_7\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNICIK32_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFJCI8_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI0VUU1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIQCIQ1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_243_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_299\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_315\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_219\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_275\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIUGIQ1_7\ : std_logic;
signal \processor_zipi8.shift_rotate_result_7\ : std_logic;
signal \processor_zipi8.spm_data_7\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNICSGN1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1211\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_0\ : std_logic;
signal \processor_zipi8.sy_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_1\ : std_logic;
signal \processor_zipi8.sy_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe23\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_123\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_99_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_5\ : std_logic;
signal \processor_zipi8.stack_memory_3\ : std_logic;
signal \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_3\ : std_logic;
signal instruction_16 : std_logic;
signal instruction_15 : std_logic;
signal \processor_zipi8.un28_carry_flag_value_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_6_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNISIMM1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe28\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI86UU1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNI2KHQ1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFG9I8_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_0_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIKPJ32_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI4QLM1_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe16\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_5_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_2_cascade_\ : std_logic;
signal instruction_7 : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.bank\ : std_logic;
signal \processor_zipi8.sy_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe29\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe27\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_4_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIKAMM1_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_271\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_311\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_295\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_1_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_215\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_239\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIASHQ1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIC2MM1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFHAI8_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIS1K32_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIGEUU1_2_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI06K32_3_cascade_\ : std_logic;
signal instruction_10 : std_logic;
signal instruction_11 : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIE0IQ1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV1BI8_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIG6MM1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIKIUU1_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_3_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe24\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe25\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_5\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_6\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe26\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_7_cascade_\ : std_logic;
signal instruction_5 : std_logic;
signal instruction_6 : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_7_cascade_\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI0NMM1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_7\ : std_logic;
signal instruction_9 : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_7\ : std_logic;
signal instruction_8 : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_3\ : std_logic;
signal \processor_zipi8.arith_logical_result_5\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5\ : std_logic;
signal \processor_zipi8.arith_logical_result_6\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_6\ : std_logic;
signal \processor_zipi8.arith_logical_result_7\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_4\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20\ : std_logic;
signal \processor_zipi8.arith_logical_result_0\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0\ : std_logic;
signal \processor_zipi8.arith_logical_result_1\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_1\ : std_logic;
signal \processor_zipi8.arith_logical_result_2\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_2\ : std_logic;
signal \processor_zipi8.arith_logical_result_3\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_3\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3\ : std_logic;
signal instruction_4 : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_3\ : std_logic;
signal \processor_zipi8.alu_mux_sel_1\ : std_logic;
signal \processor_zipi8.arith_logical_result_4\ : std_logic;
signal \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\ : std_logic;
signal \processor_zipi8.alu_mux_sel_0\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_4\ : std_logic;
signal \CLK_3P3_MHZ_c_g\ : std_logic;
signal \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_3P3_MHZ_wire\ : std_logic;
signal \LED1_wire\ : std_logic;
signal \BTN1_wire\ : std_logic;
signal \test_program.Ram2048x2_inst3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \test_program.Ram2048x2_inst0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \test_program.Ram2048x2_inst0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \CLK_3P3_MHZ_wire\ <= CLK_3P3_MHZ;
    LED1 <= \LED1_wire\;
    \BTN1_wire\ <= BTN1;
    instruction_7 <= \test_program.Ram2048x2_inst3_physical_RDATA_wire\(11);
    instruction_6 <= \test_program.Ram2048x2_inst3_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst3_physical_RADDR_wire\ <= \N__12595\&\N__12757\&\N__13003\&\N__14194\&\N__13798\&\N__14011\&\N__13648\&\N__17698\&\N__15292\&\N__15682\&\N__15505\;
    \test_program.Ram2048x2_inst3_physical_WADDR_wire\ <= \N__12592\&\N__12754\&\N__13000\&\N__14185\&\N__13795\&\N__14002\&\N__13645\&\N__17695\&\N__15277\&\N__15679\&\N__15508\;
    \test_program.Ram2048x2_inst3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \processor_zipi8.spm_data_7\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(7);
    \processor_zipi8.spm_data_6\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(6);
    \processor_zipi8.spm_data_5\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(5);
    \processor_zipi8.spm_data_4\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(4);
    \processor_zipi8.spm_data_3\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(3);
    \processor_zipi8.spm_data_2\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(2);
    \processor_zipi8.spm_data_1\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(1);
    \processor_zipi8.spm_data_0\ <= \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(0);
    \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__12197\&\N__13366\&\N__12284\&\N__19246\&\N__17186\&\N__15049\&\N__21569\&\N__16840\;
    \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__12196\&\N__13370\&\N__12283\&\N__19247\&\N__17185\&\N__15050\&\N__21565\&\N__16841\;
    \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__16701\&\N__16632\&\N__18803\&\N__21860\&\N__20056\&\N__22049\&\N__21707\&\N__21112\;
    \processor_zipi8.stack_memory_11\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(15);
    \processor_zipi8.stack_memory_10\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(14);
    \processor_zipi8.stack_memory_9\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(13);
    \processor_zipi8.stack_memory_8\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(12);
    \processor_zipi8.stack_memory_7\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(11);
    \processor_zipi8.stack_memory_6\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(10);
    \processor_zipi8.stack_memory_5\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(9);
    \processor_zipi8.stack_memory_4\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(8);
    \processor_zipi8.stack_memory_3\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(7);
    \processor_zipi8.stack_memory_2\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(6);
    \processor_zipi8.stack_memory_1\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(5);
    \processor_zipi8.stack_memory_0\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(4);
    \processor_zipi8.stack_i.stack_bit\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(3);
    \processor_zipi8.stack_i.stack_bank\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(2);
    \processor_zipi8.stack_i.stack_zero_flag\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(1);
    \processor_zipi8.stack_i.data_out_ram_0\ <= \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\(0);
    \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&\N__15779\&\N__15386\&\N__14603\&\N__13076\&\N__14690\;
    \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&\N__15166\&\N__17261\&\N__14501\&\N__14675\&\N__14582\;
    \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_WDATA_wire\ <= \N__14402\&\N__12543\&\N__12692\&\N__12944\&\N__14124\&\N__13740\&\N__13941\&\N__13596\&\N__17608\&\N__15204\&\N__15630\&\N__15450\&\N__13502\&\N__25637\&\N__18047\&\N__17992\;
    instruction_13 <= \test_program.Ram2048x2_inst6_physical_RDATA_wire\(11);
    instruction_12 <= \test_program.Ram2048x2_inst6_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst6_physical_RADDR_wire\ <= \N__12559\&\N__12721\&\N__12967\&\N__14158\&\N__13762\&\N__13975\&\N__13612\&\N__17662\&\N__15256\&\N__15646\&\N__15469\;
    \test_program.Ram2048x2_inst6_physical_WADDR_wire\ <= \N__12556\&\N__12718\&\N__12964\&\N__14149\&\N__13759\&\N__13966\&\N__13609\&\N__17659\&\N__15241\&\N__15643\&\N__15472\;
    \test_program.Ram2048x2_inst6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    instruction_3 <= \test_program.Ram2048x2_inst1_physical_RDATA_wire\(11);
    instruction_2 <= \test_program.Ram2048x2_inst1_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst1_physical_RADDR_wire\ <= \N__12619\&\N__12781\&\N__13027\&\N__14218\&\N__13822\&\N__14035\&\N__13672\&\N__17722\&\N__15314\&\N__15706\&\N__15529\;
    \test_program.Ram2048x2_inst1_physical_WADDR_wire\ <= \N__12616\&\N__12778\&\N__13024\&\N__14209\&\N__13819\&\N__14026\&\N__13669\&\N__17719\&\N__15301\&\N__15703\&\N__15532\;
    \test_program.Ram2048x2_inst1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    instruction_9 <= \test_program.Ram2048x2_inst4_physical_RDATA_wire\(11);
    instruction_8 <= \test_program.Ram2048x2_inst4_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst4_physical_RADDR_wire\ <= \N__12583\&\N__12745\&\N__12991\&\N__14182\&\N__13786\&\N__13999\&\N__13636\&\N__17686\&\N__15280\&\N__15670\&\N__15493\;
    \test_program.Ram2048x2_inst4_physical_WADDR_wire\ <= \N__12580\&\N__12742\&\N__12988\&\N__14173\&\N__13783\&\N__13990\&\N__13633\&\N__17683\&\N__15265\&\N__15667\&\N__15496\;
    \test_program.Ram2048x2_inst4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    instruction_15 <= \test_program.Ram2048x2_inst7_physical_RDATA_wire\(11);
    instruction_14 <= \test_program.Ram2048x2_inst7_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst7_physical_RADDR_wire\ <= \N__12547\&\N__12709\&\N__12955\&\N__14146\&\N__13750\&\N__13963\&\N__13600\&\N__17650\&\N__15244\&\N__15634\&\N__15457\;
    \test_program.Ram2048x2_inst7_physical_WADDR_wire\ <= \N__12544\&\N__12706\&\N__12952\&\N__14137\&\N__13747\&\N__13954\&\N__13597\&\N__17647\&\N__15228\&\N__15631\&\N__15460\;
    \test_program.Ram2048x2_inst7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    instruction_5 <= \test_program.Ram2048x2_inst2_physical_RDATA_wire\(11);
    instruction_4 <= \test_program.Ram2048x2_inst2_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst2_physical_RADDR_wire\ <= \N__12607\&\N__12769\&\N__13015\&\N__14206\&\N__13810\&\N__14023\&\N__13660\&\N__17710\&\N__15304\&\N__15694\&\N__15517\;
    \test_program.Ram2048x2_inst2_physical_WADDR_wire\ <= \N__12604\&\N__12766\&\N__13012\&\N__14197\&\N__13807\&\N__14014\&\N__13657\&\N__17707\&\N__15289\&\N__15691\&\N__15520\;
    \test_program.Ram2048x2_inst2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    instruction_17 <= \test_program.Ram2048x2_inst8_physical_RDATA_wire\(11);
    instruction_16 <= \test_program.Ram2048x2_inst8_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst8_physical_RADDR_wire\ <= \N__12536\&\N__12691\&\N__12939\&\N__14122\&\N__13729\&\N__13939\&\N__13585\&\N__17639\&\N__15234\&\N__15610\&\N__15448\;
    \test_program.Ram2048x2_inst8_physical_WADDR_wire\ <= \N__12532\&\N__12699\&\N__12951\&\N__14121\&\N__13728\&\N__13938\&\N__13584\&\N__17620\&\N__15214\&\N__15609\&\N__15437\;
    \test_program.Ram2048x2_inst8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    instruction_11 <= \test_program.Ram2048x2_inst5_physical_RDATA_wire\(11);
    instruction_10 <= \test_program.Ram2048x2_inst5_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst5_physical_RADDR_wire\ <= \N__12571\&\N__12733\&\N__12979\&\N__14170\&\N__13774\&\N__13987\&\N__13624\&\N__17674\&\N__15268\&\N__15658\&\N__15481\;
    \test_program.Ram2048x2_inst5_physical_WADDR_wire\ <= \N__12568\&\N__12730\&\N__12976\&\N__14161\&\N__13771\&\N__13978\&\N__13621\&\N__17671\&\N__15253\&\N__15655\&\N__15484\;
    \test_program.Ram2048x2_inst5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    instruction_1 <= \test_program.Ram2048x2_inst0_physical_RDATA_wire\(11);
    instruction_0 <= \test_program.Ram2048x2_inst0_physical_RDATA_wire\(3);
    \test_program.Ram2048x2_inst0_physical_RADDR_wire\ <= \N__12629\&\N__12791\&\N__13037\&\N__14225\&\N__13832\&\N__14042\&\N__13682\&\N__17732\&\N__15320\&\N__15716\&\N__15541\;
    \test_program.Ram2048x2_inst0_physical_WADDR_wire\ <= \N__12628\&\N__12790\&\N__13036\&\N__14221\&\N__13831\&\N__14038\&\N__13681\&\N__17731\&\N__15313\&\N__15715\&\N__15542\;
    \test_program.Ram2048x2_inst0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \test_program.Ram2048x2_inst0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \test_program.Ram2048x2_inst3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0010011000100001000000100010000000000010000000000000011000100100001001100000000000000000001000000000000000000001000000000000000000100000001000000010000000100000000000010000100100001000000010000000100000001000000111000001100100011000001010000001100000011001",
            INIT_E => "0000110000001100000010000000100000001001000000000001010000010100000000010000000100000101000001000000000000000000000001000000010000000100000001000000000100000100001001010000010100000100000001000000010100000000000000000000000000100110001001100000001100000011",
            INIT_D => "0000011000000110001000110010000100000000001000000010001000100000000000100000101100101000000010110001111000011111001010110000100100001000000010000010101100101001000010110000100100001010001010000010101000100000001000100010000100000000000000010010000100100001",
            INIT_C => "0010001000100010000000010000000100100001001000010000000000000000001000000010000000000000001000000010000000000000001000000001000000000000000100010010100100111000000010000001100000101000001110000000100000011001000010000011100100101000001010010001100100011001",
            INIT_B => "0001000000010000000100010000000100010001000100000000001000000010001000000010000000000000000000010001000000000001000000010000000000001000000010000001000100011000000010010000100000001000000010000000000000001000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000001000110000001000000010000000000010001000000010001000100000000000100010010000110110000000000000001000010000000000000001000000010010001100000001001000010000000100100001000000010000001100000011001000010000000100100000000000000010000000000000000",
            INIT_9 => "0000000100000000000000000000000000000000000000000000000000000001000100000001000000010010000000000001100100010000000100100000100000011000000010010001000000001000000000100000000100000100001000000001001000110000000101110011000000010010001000000000101000100000",
            INIT_8 => "0001001000110001000000100011000100100010001000000010100000100000001000000000000000100010000000100010000000000000001010010000000000001000001010000000100000101000000011010010110000001000001010000000110000101100000010010010100000000000001000000000000000100001",
            INIT_7 => "0000010000100000000100000010000000000100001000010000000000100000000000000010000000010000001000010000100000100000000000000010100000001010001110100000100000101000000000000010100100000000001001010000010000100101000011000010010100100100001001000010110000100101",
            INIT_6 => "0010010000000101001011000000010100110100000001010010010000011001000100000011010000010100001001000001010000110100000001000010010000000100001001000000010000110000000101100010001000000100001100010000010000100001000101000011100100001100001010010000100000101001",
            INIT_5 => "0000100000111000000110000010110100001100001111010000110000101000000100000011000100000010001000010000000000100101000001000011000100010000001000010000001000110111000001100010001100010100000101100000000000011010000001100000100100001000000111010001010000001101",
            INIT_4 => "0000010000010101000000000000000100010100000100010000000100010100000001010000000100000001000100000001001100000101000001000001000000000011000000000001001100010001000001000011010000000001000000100000000100110011000100000010001000000001001100100000000100100010",
            INIT_3 => "0000001000110001000100000011000000010010001100100000000100100000000000010010001000000000001000000000000100100011000010100011000000000001001100000000000000100000000100000000001000010001000100010000000000000000000000010000001100000000000000010001000000000001",
            INIT_2 => "0000000000000001000000000000000100000000000000010000000000001001000000000000000100000010000000110000100000000011000000000000000100010010000000110000000000000001000010000000000101010000000000010101001000000011011100000101000100000100000000010000000000000001",
            INIT_1 => "0000001001000011010000000000000100010000010000010001000000010001010000100100011100000000000000010000000000000001000000000100000101000010001000110000000001100001000000000010000101000000011000000000001000100010000000000010000000000000011000000100000000100000",
            INIT_0 => "0000001001100010000010000010000001000000011000000000000100100001000000100010001000000000011000000100000000000000000000010100000100000000000000000100010001000000000000000100000000000001000000000000010001000100010001000000111000000100010001000000010000000100"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst3_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst3_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst3_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst3_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst3_physical_WDATA_wire\,
            RCLKE => \N__16223\,
            RCLK => \N__33659\,
            RE => \N__22529\,
            WCLKE => \N__16222\,
            WCLK => \N__33658\,
            WE => 'L'
        );

    \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RDATA_wire\,
            RADDR => \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_RADDR_wire\,
            WADDR => \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_WADDR_wire\,
            MASK => \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_MASK_wire\,
            WDATA => \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__33619\,
            RE => \N__22562\,
            WCLKE => \N__17477\,
            WCLK => \N__33618\,
            WE => \N__22560\
        );

    \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RDATA_wire\,
            RADDR => \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_RADDR_wire\,
            WADDR => \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_WADDR_wire\,
            MASK => \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_MASK_wire\,
            WDATA => \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__33617\,
            RE => \N__22563\,
            WCLKE => \N__19070\,
            WCLK => \N__33620\,
            WE => \N__22561\
        );

    \test_program.Ram2048x2_inst6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000101000011100000011100001100100001000001111010010110000011001000010000001110100111111000111110001101000111100001111100001110100011110001111010001010000011101000111100001111100011110000111110001111000011111000010110000101100011000000111110001101000101110",
            INIT_E => "0001111000111011001110100011111100100010001001110011011000111011001010110010111000101110001010100010101000101111001011110010101100101110001010110000101100101110001011100010101000101110000010110011101000111110001010000011111100011110001110010000101100101110",
            INIT_D => "0000111000101001001010000000101100001010001011110010000000001111000011100010110000101010000010100001101000101001001011010001111000111110001111110010111100001100001011110010110000001100001011010010011100000111001001100000111000001110001011110010011100001110",
            INIT_C => "0010110000001111000001010010111000101111000011100000011000101111001011100000111000000110001011100010111000001110001101100001111000011110001111100011111100010110000111100011111100111110000111110001111000111110001111100001111000101110000111110000111100101110",
            INIT_B => "0011010000101111001011110010111000001111001011100011110000111111000111010011111100111110000111100000111000001111001111110011111000111110001101110010111100101110001101110011111000011110000111110001111000011110000111100001111000011110000111100001011000011110",
            INIT_A => "0001101000011110000101100000111100001110001111100011011000001111000011100010111000000100001011110011110000111110001111100011011100111110001111100010101000101111001111100011111000111110001111110010111000101110000111100001111100010110000111100001111000011111",
            INIT_9 => "0001111100011110000111110001111100011010000111110001111000011110001111100010111100101100001011010010111000100110001111000010110100100110001111100011110000101111001111100011110000111000001110110011111000101101001000010011101000101111001011010010101000100001",
            INIT_8 => "0010100000101001001000100010101100101010000110110011101100010011001110110001101100110000000110110010100000011011001111110001011000111110000111110010101000101011001010110010101000101010001010110010101000101011001010100010101100100110001011110010101100101110",
            INIT_7 => "0010111100101011001111100010111100111010001111110011111000111111001111100011111100101101001011100011111000110111001111100011111100110100001011110010110000111111001010100010111100101110001011110010111000101111001011100010011100101110000011110010011000001111",
            INIT_6 => "0010111000001111001011100000011100101110000011110011011000001011000010100001111100100110001000110010011000100011001001100010001100100110001100110011011000100011001001000010001100110100001000110010001000110011001010100010001100101010001010110010111000111111",
            INIT_5 => "0011101000101111001011100010101100111010001010110010101000111011001001000010111100101010001011110010111000111001001110100010111100101110001011110011110000101011001010100001100100001010001010010000110000000111000010110001110000010101000010100000100000001001",
            INIT_4 => "0001100100001000000011000001110100000001000011000000110000001000000010000001110000011100000011000000111000001000000110000000111100001110000111000000111000001100001011000000111100001010001110000011110000101110001011100010110100111100001011100010111000111100",
            INIT_3 => "0011011000100101001011000011111100101110001011000010010000101110001011100010000000100101001011100010101000100100001001100010110000111000001111100010111100111010001110100010110100110000001100100010001000110011001100100011000100110011001100010011000100100011",
            INIT_2 => "0011001101110001011000010001001100010011011100110001111100111011000111010001110100001001000111010001000100011001000110010001001100010001000010010000101100010011000100010001101100111001000010110000000100111001001110110000101100011001001110110011100101111111",
            INIT_1 => "0111100100101101001011110011101101111101001011110010100101101111001111010011100100111111001110110001100101111011010011010011111100111001001111010111111100111011001000010110011100101101001011110010110100101101001000110110111101101101001000110010000100101111",
            INIT_0 => "0110110100100101001001110110111100101100001111110011110000101110001011000111110101110110001001110010010000110111011101000010011000100100011101110010000000110011001101000011001100110110011101000111010100110010000111010011101001011101001110100001110101111010"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst6_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst6_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst6_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst6_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst6_physical_WDATA_wire\,
            RCLKE => \N__16225\,
            RCLK => \N__33694\,
            RE => \N__22556\,
            WCLKE => \N__16224\,
            WCLK => \N__33693\,
            WE => 'L'
        );

    \test_program.Ram2048x2_inst1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0010000000101000000000000000100100000000001000000010010000000110000000100000001000000001001000010000000000100010000000000010001000100000001000000010000000110000000010000011101000001000001110100000101000111000000010110010100100001000000010000000100000001010",
            INIT_E => "0000100000001010000100000000001000000000001010100000000000100000000000000010000100000100001001000000000000000000000011100000111000001110000010100000101000001010000010110000101100001011000101000000001000000000001000100000000000110100001101000000000000000011",
            INIT_D => "0000000000000000000000010000010100000010000000000010000000100000000010110000101000101010001111100000111000011011001111010010100000111110000110000000110100001000001011000000100100100001001000000010100100001101000000010010010000001010000001010000000000010100",
            INIT_C => "0000101000100010000000000000000000001001001000110000000100000010000011010000011100000101000001110010110100010101001001010011010100001100000101000010110000110100000011110000111000101110000010100000111100001010000011100010101000001110000010010000111000001100",
            INIT_B => "0010111000001100001111100001110000011111000110010001111100001010001111010010100100001101000000100000100000000011000110010010011000011000001011100010100100001100001000000000010100000001000000000001100100011001000110110001001100011011000100110001001100010011",
            INIT_A => "0001101000000010000001100010010000001111000001000010011100000000000111110001000000010111000100100010110100110000001010010001111000101001000011100010100100001010001010010001101000001000001110000000100100101000001111010001110000111101000011000011110100001110",
            INIT_9 => "0011110100001110001111000000101000101000000110100010100100110000001010000010000000111000000100000011000000010000001110000001110000100001000001000001100100111100000110010010011000011011001000010001110000100110000100000011000000011100000101000000000000011000",
            INIT_8 => "0001100000000000000100000001000000001000000000000000001000001000000110000001000000000010000000100000100000000100000011000000111000011000000110100001100000101110000110010010101000011001001011000001100000001000000110000000110100011100000011000001000100001011",
            INIT_7 => "0001000000111010000101000011111000000000001010100001000100010000000000000000000000000011000000000000000000000001001110000011100000110010001100100010000100000000001010000000101100100100000001110010010100000111000001010010111100001100000001000000010000000101",
            INIT_6 => "0000110000000101000001000001110000001000000000110001000000000011000110010001001000101000001000100011100000111000001010000000000000111000000010000011100000000000001010100000101100001001001100010011100000101000001110000011111000101100000011100011110100001110",
            INIT_5 => "0011100000001010001010010000100100001100001011010001110000101100000111000011110100000001001010010001010100001101000100000000100000000111000010010001001000000011000100000010010100010001000100100000010100000101000110100000100000010001000000010000110000001100",
            INIT_4 => "0000000000000000000101000000010000010001000100010000100000001000000110010000000100011000000000010000101000000111000110000000000000010110000010010001111000111111000010010010100000001000000110110011110000101101001011100010010000101100000100010010010100011010",
            INIT_3 => "0011011000000010001111000001100000011011001101100000000100110101000011000011110000000001001100000000100100011011000001110000011000011011000100010000010100001010001100000011101000111111000100010011111100011001001011010000001100111101000110010001110100110001",
            INIT_2 => "0001111100111000000011010100000000011111000111000000111100001100001010000000001100100010000000010011011000010011001011000000000100110100000100100010110000000000001101000111001000111100001100000000010100000011011001010110010100010001001001110111100100101000",
            INIT_1 => "0110110100001010001010010000100000111001010110100110010000001001010100000111111100000000001010010100000000001011010000000000000000110000001100100010110000100010011100000000000001111101010010010011000100000010011100010000001001010001001001010001000100100000",
            INIT_0 => "0101010100100011010100000011001001001100010001000001110000010100010011010000001001011001000101100000100000001100000111000001000001101100001010000110100001100010001110000011110001111001001100000111100000001001000110000000100101010000000000110101100000000001"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst1_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst1_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst1_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst1_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst1_physical_WDATA_wire\,
            RCLKE => \N__16231\,
            RCLK => \N__33696\,
            RE => \N__22501\,
            WCLKE => \N__16230\,
            WCLK => \N__33695\,
            WE => 'L'
        );

    \test_program.Ram2048x2_inst4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011101000000011000111100001110100101000000010110000111000010000001001110000110000000101000101000000101000101001001111110001010000010100001010110010000100010101000010110000100000011110000101100001010100001000000000010001011000011001000110010011100000010001",
            INIT_E => "0001010100001010000100100011000100001011000000100000010000000000000000000001011000000110000010000000101000010010000011010000100000000100000100110000001100001001000011100011001000001100001010010010100000011011000010100010000000100100001010100000001000000100",
            INIT_D => "0011110000111010000110000010001000100010000111000000001000100011001110000001101000011110001001110010010100001011000001100010000000001011001011110000110000100010000100100011110000110111000000010000110100110101000000000010011000110100000100010001010000100110",
            INIT_C => "0000001000100011001100000001010000010100001000000010010000010111000000100010000100010010001100110001010000100001000101000010011100110011000101010000111000101011001001000001110000011000001000100001101000111100000001100010001100000101001011010000100000110110",
            INIT_B => "0010111100001001000001100011110000001010000000100001101100111111000101010000000100010100001111000001100000000011001110100001100000111010001011110000110000011000000011000010011000001010000100010011101000101111001111000001000100001100001011110000001000010001",
            INIT_A => "0011001100100011001000000000000000010000000001100000011000100001001001100001011000100010001000110001000000010100000111000010100100110100000111100011101000100001000110100001101000010000001001010010010000011010000011100000010100001010001110100011000000001101",
            INIT_9 => "0011110000110010000011110000110100000011001100100011000000001100000011000000011000001110001110010010101100001101001010100010101000011110000001100000110000101001001110000000011000001000000111010000010000100010001101000001011000100101001101110001101100011100",
            INIT_8 => "0001001100100001001100010001010000100000000000100000100000101100000000000001001000100010001101100010000000000001000010000010110000000000000100100000001100001001000011100011001000111001000010000011010100110010000000110000100100001010001100100011000000000000",
            INIT_7 => "0011010100111010000010100000000100001011001010100010010000010101001001000011101100001010000001000000101100101000000011110001111000001110001000110010100000010101001110000011100100011100000001110000111000111001001010100000111100110000000100010001010000100111",
            INIT_6 => "0000011000010001001010100010111100100000000100010000010000100011000101100000010100110110001001110001010000001001000000000010011100110010000010010010011000100111000101100000101100000000001001010000000000011011000111000010100100100100000000010011000000101001",
            INIT_5 => "0000100000000001000111000010100100100100000001010010010000111001000110000000000100000000001000110011010000001011001010100010000100011000000010110000011000100011000001000011101100111100000001110000101000101001000110000000101000101110001000000011110000001111",
            INIT_4 => "0000110000100100000010000001101100110000001000000010010000000010000100000010100000001000000000100011110000101010001000100000000100000000001110100001000000000010000000100010100100111000000000100000111000001000000100000010011100100100000010100010110000110110",
            INIT_3 => "0000100100000010000010110011010100111100000000110010011000100100000011000000101000000000001001100010100000001010001001000010001100010110000100100001111000100010000010010000101100011010001100100011101100001110001111000010001100011100000111100000101000100000",
            INIT_2 => "0010100000001110010011000010001000101110011111000110110001001010010010100001011000000010011000000010001000010010011010000110110001000100000000000000111001101110001010000000101000001010011011000101010000010000010101100011011000110100001010100101101000010100",
            INIT_1 => "0000100000101000011101100001001000100000001011100000001001000000010001000011100000101010000001100110100000011010001001100010010001000100000110000000111000100010001010000100001001101010001100000001100000000100010100100011001000101100000010100110001000110000",
            INIT_0 => "0001100000001000000100100111001001110000000101100010111000100100010111000001110000001110001000110100110100001110000010100010000000111000010111000110110000100011000011010000101001001000001100100011111000001100011111100011100000001000000001100000000001110010"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst4_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst4_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst4_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst4_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst4_physical_WDATA_wire\,
            RCLKE => \N__16218\,
            RCLK => \N__33657\,
            RE => \N__22530\,
            WCLKE => \N__16219\,
            WCLK => \N__33660\,
            WE => 'L'
        );

    \test_program.Ram2048x2_inst7_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0010010100111001011011110111110100101100001001000010110000101100001011000010100000100110001010000011010000011000001001000000100001110100010110100010001000011010001101000001110000110000000111100011011000011100000101000001010000011110000101100101110001011100",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000101000001011000010110000101100000010000000100000000000000101000001010001010100010100000100100011000000110111000100110001000100110011001100110001001100010011000100100011100100010010001110010001001100111001000000100011100000000001000010100000001000011011",
            INIT_E => "0001001100101011001100110010101100100010001100110010001000101011001011110011111000101011001111110010111000111110001010100011100000101010001110000000111100011101000010100001100000001010001111000010011000000100001000000000011100000000000000010000000000110000",
            INIT_D => "0000010000010010000000110011011100100011001100000000000000110110001000000011110000000000001110000010000000101010000101100001111000100110001011000000010000011010001001010001100000000101000111010000010000010100000001000011110000101110001111000000011000011100",
            INIT_C => "0000110000110100001001000011111000001111001111100010011100111111000011100001011100100110001111110000111000011011000101100010101100111110001001100001011100100110001111100010110000011110000011010011111000101100000111100000110000001110000111000010111000101000",
            INIT_B => "0010110000001010001011100000000000001111001000000011110100010001001111000001001000011110000000100001111000000010001111100000001000110110000010100010111000001010001111110000101000010111001000110001011000100011000111100010000100011110001000010001001000101101",
            INIT_A => "0001101000101100000001100011100100011110001100000000011000001000000011100000100000000100000010000011110000110010001101100011101000111110001010100011101000101110001111100010101000111110001010100010111000101010000111100010101000011110001010100001111000100000",
            INIT_9 => "0001111000100000000111100010000000011010001001000001111000100100001011100000010000101101000001110010011000001101001011000001111100111110000111000010010000010100001111000000010000111000001001000010110000101001001100100011111100101001001000100010000100100100",
            INIT_8 => "0010100000101100001000000010110000001000000101010001001100010100000110110001110000000000000011010000100100000110000101100000001000011110000010100010101100011010001010100001101100101011000110110010101100011010001010100001101000101110000111110010101000010001",
            INIT_7 => "0010101100010000001011110000010000111010000100000011101000010000001110110000000100111000000000110011001100001001001110110010100000101000001110000011000000100010001000100011001000101010001101100010101000110110001000100011011000001010000111100000001000011110",
            INIT_6 => "0000101000010110000000100001011000001010000011000000001000001000000111100001010000100010000010000010001000001000001000100000100000100010000010000010001000001000001000000000100000100000000010100011001000111010001000100010101000101010001010100010111000101110",
            INIT_5 => "0010101000101010001010100010101000101010001010100011101000111010001011000010110000101000001000000010100000100000001011100010010000101110001000000010100000100000000110000011000000101000000000100000011000101110000010000010101000001010001010110000000100100011",
            INIT_4 => "0000100000100010000111010011011100000000001010100000100000101010000011000010111000001100001010100000100000101010000011100010111000011100001110000000110000100110000010100000001000101000001001100010111000000010001011000000010000101110000001100011110000011100",
            INIT_3 => "0010010000001110001101100001011000101100000001100010011000010110001000000001010000100110000100100010010000011000001011000000110000101010000000100010101000001001001011010010110100110010001111100011001000111100001100000010110000110001001011110010001100101111",
            INIT_2 => "0011000101111101000000110100111101010011000111010001001101010001000011010110000100001101011010010001000101100101000100010110011100000001011101010001001101111101000110010110110100001001001001010011000100111101000010110000110100111001001010010011100100001001",
            INIT_1 => "0010100100001001001111110001100100101101000011010110110101010101001110010001000100111111000100010000110100000001000010010000000100111001001000010011101100101101011001010111110100100101001100010010100100110001001000110011000100100001001101010010010100110101"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst7_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst7_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst7_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst7_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst7_physical_WDATA_wire\,
            RCLKE => \N__16229\,
            RCLK => \N__33707\,
            RE => \N__22567\,
            WCLKE => \N__16228\,
            WCLK => \N__33706\,
            WE => 'L'
        );

    \test_program.Ram2048x2_inst2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000101000100011000010100010000000000000000000100010011000000100000000000010001000000001000100010000000000010001001000000001000000100010001100100000101000110000000010100001100000001010000110000000100000011010000110010001101100101000000010000001100000001011",
            INIT_E => "0001110000001110000010000011001000001000001000100001010000110110000010010010001000001100001000110000110000100010000001000010100000000100001010000000000000001000000001010000110000100100000010000010000000000000000000000010000000100010001001000000001000000010",
            INIT_D => "0000011000000000001000010000000100000000000000000000100000000000001010010000101100101111001010110001110000101111001011000010110100001101000011010010110000001101000011000000110100101100001000100000000000101000000000010010000100001000001010010010000000000001",
            INIT_C => "0000101100101011000000000010000100001000001010100010100000000010000011000010101000000000000000100000110000001010001000000010101000001000001010110000000000000011001010000000100000001000000010000010100100001001001010010010100100001000000010010001100000101000",
            INIT_B => "0010000100100001001100000010000000010001000100010000001000010010001000000011000000100001001000110011010000000011001000010001001100100001000100110001100100111011000110010010101100011000000010100000100000011010000000000001000000000000000100000000000000010000",
            INIT_A => "0000100000011001000001000000000000001101000010010000010000100000000111010000100100010110000100110011110100001001001111000000001100101101000010110011100000001010001111010000101100111101000010110011110100011011000110000000111100010001000001110001000000000101",
            INIT_9 => "0001000000000101000100000000010000010000000000000001000100000101001000000000010000110000000001000011100100011100001010100001110000101001000011010011100000001100001100010001011100010100000100000001110000011010000100000001000100011000000110000001000000001000",
            INIT_8 => "0001100000011011000010010000000000001000001010000001000000011000001110010010100100100010000010100000100000101000000101000001001000111100001011100000100000101010000011000010101000001000001010100000110000101010000010010010101000000100001000100000000100100001",
            INIT_7 => "0000000000000000000001000000000000010000000100000001000000000001000000000000000000010001000000010001000000011000000110000000100000011010000010100000100100001000000011010000101000000101000001100000010100000110000001000000111000001101001011100000010100000110",
            INIT_6 => "0010110100101111001001010000111000011101001010000001000000010000001110010011100000000101000101000000010100010000000000010001010000000001000000000001010100000100000001110001001100010000000001000000000000100011000011000011001100011000001011100000110000101010",
            INIT_5 => "0001100100101010000011010011101000011101001010110000100100101110000001010011000000010001001100000000001100100100000100110010000000000001001100100000011100110010000001100000001100000010000101000000110000001000000010100000100000011110000010000000110100011001",
            INIT_4 => "0000000000010100000001000000000100000000000100000000100000010100000010010000000100011100000000010000101000010110000010000000001100001010000001010000011000010010001101000000001000000100000000110001010000100000000001000011000000000100001000010000111000100001",
            INIT_3 => "0001011000100011000101000011001000000100001100000000011000100000000011010010100000000011001010010000101100101011000101100011001000011100001110000000111100100101001011100000001000110001000100000010000000000010001100110001001100110010000000110010000000000011",
            INIT_2 => "0011001000010011011000000000001100010010000000110001111000011111000000100000000100001010000000110001000000000001000110000001000100000010000000110000100000000011000100000001001101100000000000010000001001000010001110000100001000111100001100100011000000011000",
            INIT_1 => "0111011000011110001001000101101001100000000010100011010000010100001100100100001000110100010101100000010000000010010000000000000000010010011000100101000000111110000000000010001000000101011001010100001100100011000000010010001101000001001011100000000101101001",
            INIT_0 => "0000011101101110000001010010011000001100011010100100010101101000000100100010111001000100001000100011010001000010001000010101010000010000001001000000010001100100000100000010000000010000001000000101010000100100000111000100100000010000000001000001000000001000"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst2_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst2_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst2_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst2_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst2_physical_WDATA_wire\,
            RCLKE => \N__16227\,
            RCLK => \N__33676\,
            RE => \N__22502\,
            WCLKE => \N__16226\,
            WCLK => \N__33675\,
            WE => 'L'
        );

    \test_program.Ram2048x2_inst8_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0110101101011000001001010101000001100100000000000011110100000000001010100100000001110000000110000000000001001000010100010101100000000010010010000101011000001000000101000000110000010111010011100101000100001110000100010100010001010011010001000001100101000100",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0010100000000010000011010000001000000000001010100010011100001100000100110010100000110010001010100001011000101010001100110010111000010001000011100011000100001110000100000010010000010001001001000001000100100100000000000010010000000010000000000000001000000000",
            INIT_E => "0010011100000000001000110000000000101010000000000010111100000100001010110001000100101110000101010010101000010001001011000001000100101100000101010000100100010000000011010001000000001100000101010000000000011000000001010001100000000111000010000010000100011100",
            INIT_D => "0000011100011111001000000011110000000000000110010010010000111001000001110001010000100100001100000001011000010011001001010000000000100100000000010000000100010000000000010001000100000100000100010010110000010000001011010011000000001100000100010010010100010000",
            INIT_C => "0010010000110001000011110001000000101111001100010000011000010001001001100011000100001110000100010010101000010001001000100010000100000110000000000010111000101000000001000000000000100101001000000000010100000000001001000000000000110100001000010001000100000000",
            INIT_B => "0001000000000001000100010000000000110001000000010001000000100001000100100010000000000011001100000000001000110001000000110000000000001010000010010001001100001000000000110000100100000010001000010000001000100001000000000010000100000000001000010000110000100101",
            INIT_A => "0000110000100000000100010011000000100001000000000011100000000000000110010000000000010000001000000011001100000000001110100000100000100011000100000010011000010000001000110000000000100010000000000011001100000000000000100010000000000011001000000000000000100000",
            INIT_9 => "0000000100100000000000000010000100000100001000010000010100100000000101010000000100010100000000010001110100001000000101010001000000000101000000000001010000010000000001110000000000100000000000000011101100010010001000010001000100110000000000010011100000000101",
            INIT_8 => "0011100000000100001100000000010000010001001001000001100100100100000110010010010000000001001101000000001000110100000010110010100000000011001000010000011000010001000001110001000100000110000100000000011000010000000001100001000000000111000100000000000100010001",
            INIT_7 => "0000010000010001000101000000000100010000000000000001000000000100000000010001010000000001000101010000100000001100001000000000110000110001000111000010001100010100001000110001010000100011000100000010001100010000001010110001000000001011001100000000001100110000",
            INIT_6 => "0000001100110000000010110011000000001001001000000001010100110100000000010010000000000001000111000001000100001100000000010000110000000001000111000001000100001100000000010001110000010011000111000010001100011100001111110000100000100111000000000010011100010000",
            INIT_5 => "0011001100000000001001110001000000110111000100000010011100010000001101010000000000100001000000000010010100010100001100010000000000100001000100000011010100010000001001110011000000010111001000100000110100101000000000110011001000010101001000010000010000110011",
            INIT_4 => "0001010100110011000001000011001100011001001000110000110100100110000010010011001000011001001000100000111100110110000110000011000000001011001100000001011100100010001000000010000000000011001100100001000100000000000001100001001000010101000100000000111100010000",
            INIT_3 => "0001011000010010000001000000000000010111000000100000010100010000000011110001011000000001000101000000101100011100000001110000001000000001000000000000110100000101001110100001001000100001000011000010000000001100001000100000110000100011000011100011000100001100",
            INIT_2 => "0111001100001110011000010100110000010001011011000001010101100100000000110111010000001011011101000000001101100100000010110110010000010011011101000000100101101100000000010110010000110001001101000000101101000100011010010010010000001101001000000000100101000000",
            INIT_1 => "0101101100010000000011010100010001011001010001000000000101000100010101110000010000010001000001000000000101010100010000010001010000100011010001000110110101000100001000010101000001100001000100000010001100010100001000010101010001101101000101000010000101010000"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst8_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst8_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst8_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst8_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst8_physical_WDATA_wire\,
            RCLKE => \N__16217\,
            RCLK => \N__33629\,
            RE => \N__22568\,
            WCLKE => \N__16216\,
            WCLK => \N__33628\,
            WE => 'L'
        );

    \test_program.Ram2048x2_inst5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0001100000001001001110000000100100111000000110010001100000111000001010000000110100001000001011010011100000000001000010000011010100101000000101010000100000010101001010000001110100101000000010000010100000001001001010000000100100111100000100010011100000010001",
            INIT_E => "0001100000010001000111000001000100010000000000010000000000000010000000000000001000000001000000100000000100000010000000000000000100000000000010010000000000001001000000000000100000000001000010100000000100001010000000000000101000110000001010000001010000001010",
            INIT_D => "0010000000110000000001110011000000000101000100100000000100010010000000000000100000000000000010110000000000011001000100100000110000110000001001110011001000100100001000100011010000100010001101010000001000110101000001100011000000000110000000010000011000100000",
            INIT_C => "0001011000100111000001000001010000000100001101000000010000010101000001000011000100000000000000010000000000000111000000000000011100000000000000110000000000010011000010010001000000001000001101000000100000010100000110000000110100001000001011110000110000011010",
            INIT_B => "0000110000011011000011000001001000001100000101100001111000010111000111000001110100011100000111000001110000011001000110000001100000010000000100010000000000011010000000000000101000100000000011110000000000101111000000000010110100000000001111010000000000110001",
            INIT_A => "0000000000010001000001000001001000000100000000100000010000110011001001000011001000100110001101110001010000010100000101000001010100011100000101000001100000010001000110000011000000011000001110110000100000111010000010000000101100001000000011100000100000000101",
            INIT_9 => "0000100000000100000010010011010000001001001110000000110000111010000010000001111000001000000111110000000100010110000000000001111000000000001010100000001000111001000000000010100000000110000010010000010000010000000100100001010000000010000101010000011000100001",
            INIT_8 => "0000011000100001000001100010000100000110001000000001011000100000000101100010000000010110000000100001010000000001000101000000000000010100000000000000000000000101000000000000000000000000000001110000000000001011000000000011111100000100001110100000010000110000",
            INIT_7 => "0000000000110001001001000001000100110100000000010011000000001111001100000000111100110000001011100011000000100111000100000000101100000010000110110001000000001001000000000001100100000000001111010000000000111101000000000011010100000000001001110000000000100011",
            INIT_6 => "0000000000100011000000000000001100010000000000010000000000010001000100000000010100011000001001010010100000000111001110000000011100111000000001110010100000010011001110100010001100101000001100010001100000000001000000000000000100010000000000010001000000000001",
            INIT_5 => "0000000000110001000100000010000100000000001110010001000000101001001000000000100100110000000000010011000000000001001000000001000100110000001000010010001000111011000100000010100100100000001010010011000000100001001100000010100000100000000110000011001000001001",
            INIT_4 => "0010001000011000001100100000100100000010001000000001001000100000000100100010000000000010001100000001000000000000000000010001100000010000000010000000010000000000000101010010000000110100001000000000000000010000000101010000100000000100000110000001010000001000",
            INIT_3 => "0000010100111100000101010010110000000100001011000001010000100101001100000000000000110000000000000011000000000000001100000000000000100000001100010011000000101000000001000001100100010100000010000001010000001001000101000000100100010100001010000000010000111100",
            INIT_2 => "0001010000101100000101000110110001110100001011000011000001101000000100000100100000010000010000000001010001000000000101000000000000000100001100000001010000100010000101000010111001000100001111100101010000010100000101000011011001110000001100100101000000010010",
            INIT_1 => "0000000001010000010000000001101000000000010110100100000000100010000100000010000001010000001000100111000000100010001100000110101001010000000010000001000001001010010000000000111000000000000011100100000000101000010000000010001000000000011100100100000000110110",
            INIT_0 => "0010000001010100011000000001001000110000000100100110010000011110011101010011110000100000011110110100000000001011000000000101101001000001000110000000000000001011010100000010101101010000001010000001000001101110010100000010111000110000010111100111000000010110"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst5_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst5_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst5_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst5_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst5_physical_WDATA_wire\,
            RCLKE => \N__16221\,
            RCLK => \N__33674\,
            RE => \N__22555\,
            WCLKE => \N__16220\,
            WCLK => \N__33673\,
            WE => 'L'
        );

    \test_program.Ram2048x2_inst0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000100000101000000010000000000000000000000000000010011000100110000000110000000000000001000000110000001000010010000100110000000000110000001100010000000100100001001010000011101000111000001010000011101100111000001010010010101100001001000010000000101000101010",
            INIT_E => "0001111100011000000000000000011100101000001010000010001000000010000010100010010100000000000011100010000000100001001010100000111000001010001001010000000000001010000000000000000100011110000010100010001000100000000000000001000000110110001100100000001100000110",
            INIT_D => "0000011000000000000001010010010100000000000000110010000000100001000010000000101000011010000010100000110100001001000011010000100000011100000111000000110000001101000011010000100100100101001000000000110100100101000001000000000000001001000011010001000100101000",
            INIT_C => "0000111000001110000001000000000100001011000011110000001100000000000010010010111000000101000001000011101100001110000101110000010000001100000110100010100000101100000110100001101000111110000011000000110000011010001010000010110000101011001010110000111100011000",
            INIT_B => "0011100000101100001110000000101100001101000001010010011100111010001100010010010100001010000010100000111100000001000001010011111000011100000010000010101000001111000000110011000100000101000001100001110100011000000100110000111000000011000100000000000100000110",
            INIT_A => "0001100000011000001000100000011000001010000010000011010000000110000111000010100000000011001001110000100000001000001001110011111100101110000010000000100100101010000011000000100000101011001111100010101000001000000011010000111100011100000110000001101100001111",
            INIT_9 => "0000101000010001000001000000111000010000000100010011101000001010000110100000010000110100001010000010010000001110000010000010100000000000000001000010110100111000001101100001111000110000000000010001111000110000000100000001100000111100001001000010000000000001",
            INIT_8 => "0001100000100001000100000000000000001000000000000000000000000001000110000001000100000010000000100000110000010001000001110000111100011010000110000010110000001111000011000010110100001110000011100010111000101100001011010000111100001100001010000000101100001010",
            INIT_7 => "0011111000000000000001000011101100000000000000010011101000111011001010100000000000000000001010000000000000001010000110000011100000010010000000100010000000110001001010100000101100000110001011000000010100000111001001000010010100001110000001100000011100000101",
            INIT_6 => "0000110000000111000101010000010000001010000000110000001000000000000110000001001000000000001000000000101000010011001000100010000100101000000000110001000000110000000010110000001000110000001100010000100100100001000011100001111000101111001010010010110100001011",
            INIT_5 => "0001100000111000000011110000111100101010001011000010110000001010000011000011100100001000000010010010110100100101001100110001101100000000001000000000111000011111001011110000010100000101001111100000110000001001000010110000100000010100000101000000100100001101",
            INIT_4 => "0001010100001100000001010000000100000000000100000000010100000000000010000000100100011100000101000000010000001101000100000001000000001010000010000010100000011101000010000000000000000010000010000001000000110101000010000000100000101100001001000010110000000011",
            INIT_3 => "0001000100110101000110000001100000100110001111100011010100010000000100000011111000010001000100000011001000110111001000000000010000011001001110000000001100011101000000100001001100110000001100010011101100010011000000100010001000011010000100110010000000110000",
            INIT_2 => "0010101100000001000000010111000000011110011100110000101000101000000000010000100100001011000111000001001000010001000010000000000000000001000100110000000100011000011000100000001100100000001100000000000100100010000001000110101100010110001101000001100100001001",
            INIT_1 => "0110100101110010001000100000110101000000011100100000100100001001001111010111011000100010000010110000000000000000010010010101100100011001001101100000100000001101001000100010011000101100010011000000000100101011000000010000011001101011011010000010000000000101",
            INIT_0 => "0000110001100011000100110000000000101100011001100011110100000001000000000010101001000010010101100000100000100000010101010000000100101000001001000010000001000000000011000011010000000011000000110111100001110010000110000000100001000000010110000000000000000010"
        )
    port map (
            RDATA => \test_program.Ram2048x2_inst0_physical_RDATA_wire\,
            RADDR => \test_program.Ram2048x2_inst0_physical_RADDR_wire\,
            WADDR => \test_program.Ram2048x2_inst0_physical_WADDR_wire\,
            MASK => \test_program.Ram2048x2_inst0_physical_MASK_wire\,
            WDATA => \test_program.Ram2048x2_inst0_physical_WDATA_wire\,
            RCLKE => \N__16233\,
            RCLK => \N__33709\,
            RE => \N__22479\,
            WCLKE => \N__16232\,
            WCLK => \N__33708\,
            WE => 'L'
        );

    \CLK_3P3_MHZ_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__39684\,
            GLOBALBUFFEROUTPUT => \CLK_3P3_MHZ_c_g\
        );

    \CLK_3P3_MHZ_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39686\,
            DIN => \N__39685\,
            DOUT => \N__39684\,
            PACKAGEPIN => \CLK_3P3_MHZ_wire\
        );

    \CLK_3P3_MHZ_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39686\,
            PADOUT => \N__39685\,
            PADIN => \N__39684\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39675\,
            DIN => \N__39674\,
            DOUT => \N__39673\,
            PACKAGEPIN => \LED1_wire\
        );

    \LED1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39675\,
            PADOUT => \N__39674\,
            PADIN => \N__39673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21032\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BTN1_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39666\,
            DIN => \N__39665\,
            DOUT => \N__39664\,
            PACKAGEPIN => \BTN1_wire\
        );

    \BTN1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39666\,
            PADOUT => \N__39665\,
            PADIN => \N__39664\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BTN1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__10148\ : CascadeMux
    port map (
            O => \N__39647\,
            I => \N__39639\
        );

    \I__10147\ : CascadeMux
    port map (
            O => \N__39646\,
            I => \N__39632\
        );

    \I__10146\ : CascadeMux
    port map (
            O => \N__39645\,
            I => \N__39627\
        );

    \I__10145\ : CascadeMux
    port map (
            O => \N__39644\,
            I => \N__39623\
        );

    \I__10144\ : CascadeMux
    port map (
            O => \N__39643\,
            I => \N__39620\
        );

    \I__10143\ : CascadeMux
    port map (
            O => \N__39642\,
            I => \N__39616\
        );

    \I__10142\ : InMux
    port map (
            O => \N__39639\,
            I => \N__39613\
        );

    \I__10141\ : CascadeMux
    port map (
            O => \N__39638\,
            I => \N__39610\
        );

    \I__10140\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39605\
        );

    \I__10139\ : CascadeMux
    port map (
            O => \N__39636\,
            I => \N__39602\
        );

    \I__10138\ : CascadeMux
    port map (
            O => \N__39635\,
            I => \N__39599\
        );

    \I__10137\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39588\
        );

    \I__10136\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39585\
        );

    \I__10135\ : InMux
    port map (
            O => \N__39630\,
            I => \N__39582\
        );

    \I__10134\ : InMux
    port map (
            O => \N__39627\,
            I => \N__39579\
        );

    \I__10133\ : InMux
    port map (
            O => \N__39626\,
            I => \N__39576\
        );

    \I__10132\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39572\
        );

    \I__10131\ : InMux
    port map (
            O => \N__39620\,
            I => \N__39569\
        );

    \I__10130\ : CascadeMux
    port map (
            O => \N__39619\,
            I => \N__39565\
        );

    \I__10129\ : InMux
    port map (
            O => \N__39616\,
            I => \N__39562\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__39613\,
            I => \N__39559\
        );

    \I__10127\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39556\
        );

    \I__10126\ : InMux
    port map (
            O => \N__39609\,
            I => \N__39553\
        );

    \I__10125\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39550\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__39605\,
            I => \N__39547\
        );

    \I__10123\ : InMux
    port map (
            O => \N__39602\,
            I => \N__39539\
        );

    \I__10122\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39536\
        );

    \I__10121\ : CascadeMux
    port map (
            O => \N__39598\,
            I => \N__39532\
        );

    \I__10120\ : CascadeMux
    port map (
            O => \N__39597\,
            I => \N__39529\
        );

    \I__10119\ : InMux
    port map (
            O => \N__39596\,
            I => \N__39526\
        );

    \I__10118\ : InMux
    port map (
            O => \N__39595\,
            I => \N__39523\
        );

    \I__10117\ : CascadeMux
    port map (
            O => \N__39594\,
            I => \N__39520\
        );

    \I__10116\ : CascadeMux
    port map (
            O => \N__39593\,
            I => \N__39517\
        );

    \I__10115\ : InMux
    port map (
            O => \N__39592\,
            I => \N__39514\
        );

    \I__10114\ : InMux
    port map (
            O => \N__39591\,
            I => \N__39511\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__39588\,
            I => \N__39508\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__39585\,
            I => \N__39503\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__39582\,
            I => \N__39503\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__39579\,
            I => \N__39498\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__39576\,
            I => \N__39498\
        );

    \I__10108\ : CascadeMux
    port map (
            O => \N__39575\,
            I => \N__39495\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__39572\,
            I => \N__39489\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__39569\,
            I => \N__39489\
        );

    \I__10105\ : InMux
    port map (
            O => \N__39568\,
            I => \N__39486\
        );

    \I__10104\ : InMux
    port map (
            O => \N__39565\,
            I => \N__39483\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__39562\,
            I => \N__39478\
        );

    \I__10102\ : Span4Mux_v
    port map (
            O => \N__39559\,
            I => \N__39478\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__39556\,
            I => \N__39469\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__39553\,
            I => \N__39469\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__39550\,
            I => \N__39469\
        );

    \I__10098\ : Span4Mux_v
    port map (
            O => \N__39547\,
            I => \N__39469\
        );

    \I__10097\ : CascadeMux
    port map (
            O => \N__39546\,
            I => \N__39466\
        );

    \I__10096\ : InMux
    port map (
            O => \N__39545\,
            I => \N__39463\
        );

    \I__10095\ : InMux
    port map (
            O => \N__39544\,
            I => \N__39460\
        );

    \I__10094\ : CascadeMux
    port map (
            O => \N__39543\,
            I => \N__39457\
        );

    \I__10093\ : CascadeMux
    port map (
            O => \N__39542\,
            I => \N__39454\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__39539\,
            I => \N__39451\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__39536\,
            I => \N__39447\
        );

    \I__10090\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39444\
        );

    \I__10089\ : InMux
    port map (
            O => \N__39532\,
            I => \N__39441\
        );

    \I__10088\ : InMux
    port map (
            O => \N__39529\,
            I => \N__39438\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__39526\,
            I => \N__39435\
        );

    \I__10086\ : LocalMux
    port map (
            O => \N__39523\,
            I => \N__39432\
        );

    \I__10085\ : InMux
    port map (
            O => \N__39520\,
            I => \N__39429\
        );

    \I__10084\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39426\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__39514\,
            I => \N__39423\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__39511\,
            I => \N__39416\
        );

    \I__10081\ : Span4Mux_s3_h
    port map (
            O => \N__39508\,
            I => \N__39416\
        );

    \I__10080\ : Span4Mux_v
    port map (
            O => \N__39503\,
            I => \N__39416\
        );

    \I__10079\ : Span4Mux_s3_v
    port map (
            O => \N__39498\,
            I => \N__39413\
        );

    \I__10078\ : InMux
    port map (
            O => \N__39495\,
            I => \N__39410\
        );

    \I__10077\ : InMux
    port map (
            O => \N__39494\,
            I => \N__39407\
        );

    \I__10076\ : Span4Mux_s3_v
    port map (
            O => \N__39489\,
            I => \N__39402\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__39486\,
            I => \N__39402\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__39483\,
            I => \N__39395\
        );

    \I__10073\ : Span4Mux_s0_h
    port map (
            O => \N__39478\,
            I => \N__39395\
        );

    \I__10072\ : Span4Mux_v
    port map (
            O => \N__39469\,
            I => \N__39395\
        );

    \I__10071\ : InMux
    port map (
            O => \N__39466\,
            I => \N__39392\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__39463\,
            I => \N__39389\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__39460\,
            I => \N__39386\
        );

    \I__10068\ : InMux
    port map (
            O => \N__39457\,
            I => \N__39383\
        );

    \I__10067\ : InMux
    port map (
            O => \N__39454\,
            I => \N__39380\
        );

    \I__10066\ : Span4Mux_v
    port map (
            O => \N__39451\,
            I => \N__39377\
        );

    \I__10065\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39374\
        );

    \I__10064\ : Sp12to4
    port map (
            O => \N__39447\,
            I => \N__39369\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__39444\,
            I => \N__39369\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__39441\,
            I => \N__39366\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__39438\,
            I => \N__39359\
        );

    \I__10060\ : Span4Mux_v
    port map (
            O => \N__39435\,
            I => \N__39359\
        );

    \I__10059\ : Span4Mux_h
    port map (
            O => \N__39432\,
            I => \N__39359\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__39429\,
            I => \N__39350\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__39426\,
            I => \N__39350\
        );

    \I__10056\ : Span4Mux_h
    port map (
            O => \N__39423\,
            I => \N__39350\
        );

    \I__10055\ : Span4Mux_h
    port map (
            O => \N__39416\,
            I => \N__39350\
        );

    \I__10054\ : Span4Mux_h
    port map (
            O => \N__39413\,
            I => \N__39345\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__39410\,
            I => \N__39345\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__39407\,
            I => \N__39342\
        );

    \I__10051\ : Span4Mux_v
    port map (
            O => \N__39402\,
            I => \N__39335\
        );

    \I__10050\ : Span4Mux_h
    port map (
            O => \N__39395\,
            I => \N__39335\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__39392\,
            I => \N__39335\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__39389\,
            I => \N__39330\
        );

    \I__10047\ : Span4Mux_v
    port map (
            O => \N__39386\,
            I => \N__39330\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__39383\,
            I => \N__39321\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__39380\,
            I => \N__39321\
        );

    \I__10044\ : Sp12to4
    port map (
            O => \N__39377\,
            I => \N__39321\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__39374\,
            I => \N__39321\
        );

    \I__10042\ : Span12Mux_s5_v
    port map (
            O => \N__39369\,
            I => \N__39318\
        );

    \I__10041\ : Span4Mux_s3_h
    port map (
            O => \N__39366\,
            I => \N__39313\
        );

    \I__10040\ : Span4Mux_h
    port map (
            O => \N__39359\,
            I => \N__39313\
        );

    \I__10039\ : Span4Mux_v
    port map (
            O => \N__39350\,
            I => \N__39308\
        );

    \I__10038\ : Span4Mux_s3_v
    port map (
            O => \N__39345\,
            I => \N__39308\
        );

    \I__10037\ : Span4Mux_h
    port map (
            O => \N__39342\,
            I => \N__39303\
        );

    \I__10036\ : Span4Mux_h
    port map (
            O => \N__39335\,
            I => \N__39303\
        );

    \I__10035\ : Odrv4
    port map (
            O => \N__39330\,
            I => \processor_zipi8.arith_logical_result_1\
        );

    \I__10034\ : Odrv12
    port map (
            O => \N__39321\,
            I => \processor_zipi8.arith_logical_result_1\
        );

    \I__10033\ : Odrv12
    port map (
            O => \N__39318\,
            I => \processor_zipi8.arith_logical_result_1\
        );

    \I__10032\ : Odrv4
    port map (
            O => \N__39313\,
            I => \processor_zipi8.arith_logical_result_1\
        );

    \I__10031\ : Odrv4
    port map (
            O => \N__39308\,
            I => \processor_zipi8.arith_logical_result_1\
        );

    \I__10030\ : Odrv4
    port map (
            O => \N__39303\,
            I => \processor_zipi8.arith_logical_result_1\
        );

    \I__10029\ : CascadeMux
    port map (
            O => \N__39290\,
            I => \N__39286\
        );

    \I__10028\ : CascadeMux
    port map (
            O => \N__39289\,
            I => \N__39279\
        );

    \I__10027\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39276\
        );

    \I__10026\ : CascadeMux
    port map (
            O => \N__39285\,
            I => \N__39273\
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__39284\,
            I => \N__39270\
        );

    \I__10024\ : CascadeMux
    port map (
            O => \N__39283\,
            I => \N__39267\
        );

    \I__10023\ : CascadeMux
    port map (
            O => \N__39282\,
            I => \N__39264\
        );

    \I__10022\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39255\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__39276\,
            I => \N__39252\
        );

    \I__10020\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39249\
        );

    \I__10019\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39244\
        );

    \I__10018\ : InMux
    port map (
            O => \N__39267\,
            I => \N__39237\
        );

    \I__10017\ : InMux
    port map (
            O => \N__39264\,
            I => \N__39234\
        );

    \I__10016\ : InMux
    port map (
            O => \N__39263\,
            I => \N__39230\
        );

    \I__10015\ : CascadeMux
    port map (
            O => \N__39262\,
            I => \N__39221\
        );

    \I__10014\ : InMux
    port map (
            O => \N__39261\,
            I => \N__39218\
        );

    \I__10013\ : CascadeMux
    port map (
            O => \N__39260\,
            I => \N__39215\
        );

    \I__10012\ : InMux
    port map (
            O => \N__39259\,
            I => \N__39212\
        );

    \I__10011\ : InMux
    port map (
            O => \N__39258\,
            I => \N__39209\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__39255\,
            I => \N__39202\
        );

    \I__10009\ : Span4Mux_h
    port map (
            O => \N__39252\,
            I => \N__39202\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__39249\,
            I => \N__39202\
        );

    \I__10007\ : CascadeMux
    port map (
            O => \N__39248\,
            I => \N__39199\
        );

    \I__10006\ : InMux
    port map (
            O => \N__39247\,
            I => \N__39195\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__39244\,
            I => \N__39192\
        );

    \I__10004\ : InMux
    port map (
            O => \N__39243\,
            I => \N__39189\
        );

    \I__10003\ : InMux
    port map (
            O => \N__39242\,
            I => \N__39185\
        );

    \I__10002\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39182\
        );

    \I__10001\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39179\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__39237\,
            I => \N__39172\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__39234\,
            I => \N__39172\
        );

    \I__9998\ : CascadeMux
    port map (
            O => \N__39233\,
            I => \N__39169\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__39230\,
            I => \N__39166\
        );

    \I__9996\ : CascadeMux
    port map (
            O => \N__39229\,
            I => \N__39163\
        );

    \I__9995\ : CascadeMux
    port map (
            O => \N__39228\,
            I => \N__39160\
        );

    \I__9994\ : CascadeMux
    port map (
            O => \N__39227\,
            I => \N__39157\
        );

    \I__9993\ : InMux
    port map (
            O => \N__39226\,
            I => \N__39154\
        );

    \I__9992\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39151\
        );

    \I__9991\ : InMux
    port map (
            O => \N__39224\,
            I => \N__39148\
        );

    \I__9990\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39145\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__39218\,
            I => \N__39142\
        );

    \I__9988\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39139\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__39212\,
            I => \N__39136\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__39209\,
            I => \N__39131\
        );

    \I__9985\ : Span4Mux_s2_h
    port map (
            O => \N__39202\,
            I => \N__39131\
        );

    \I__9984\ : InMux
    port map (
            O => \N__39199\,
            I => \N__39128\
        );

    \I__9983\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39124\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39121\
        );

    \I__9981\ : Span4Mux_v
    port map (
            O => \N__39192\,
            I => \N__39116\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__39189\,
            I => \N__39116\
        );

    \I__9979\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39113\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__39185\,
            I => \N__39110\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__39182\,
            I => \N__39107\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__39179\,
            I => \N__39104\
        );

    \I__9975\ : InMux
    port map (
            O => \N__39178\,
            I => \N__39101\
        );

    \I__9974\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39098\
        );

    \I__9973\ : Span4Mux_h
    port map (
            O => \N__39172\,
            I => \N__39095\
        );

    \I__9972\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39091\
        );

    \I__9971\ : IoSpan4Mux
    port map (
            O => \N__39166\,
            I => \N__39088\
        );

    \I__9970\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39085\
        );

    \I__9969\ : InMux
    port map (
            O => \N__39160\,
            I => \N__39082\
        );

    \I__9968\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39079\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__39154\,
            I => \N__39074\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__39151\,
            I => \N__39074\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__39148\,
            I => \N__39071\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__39145\,
            I => \N__39068\
        );

    \I__9963\ : Span4Mux_s2_h
    port map (
            O => \N__39142\,
            I => \N__39059\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__39139\,
            I => \N__39059\
        );

    \I__9961\ : Span4Mux_s2_h
    port map (
            O => \N__39136\,
            I => \N__39059\
        );

    \I__9960\ : Span4Mux_v
    port map (
            O => \N__39131\,
            I => \N__39059\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__39128\,
            I => \N__39056\
        );

    \I__9958\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39053\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__39124\,
            I => \N__39049\
        );

    \I__9956\ : Span4Mux_h
    port map (
            O => \N__39121\,
            I => \N__39044\
        );

    \I__9955\ : Span4Mux_s1_h
    port map (
            O => \N__39116\,
            I => \N__39044\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__39113\,
            I => \N__39039\
        );

    \I__9953\ : Span4Mux_s1_h
    port map (
            O => \N__39110\,
            I => \N__39039\
        );

    \I__9952\ : Span4Mux_h
    port map (
            O => \N__39107\,
            I => \N__39032\
        );

    \I__9951\ : Span4Mux_h
    port map (
            O => \N__39104\,
            I => \N__39032\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__39101\,
            I => \N__39032\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__39098\,
            I => \N__39029\
        );

    \I__9948\ : Sp12to4
    port map (
            O => \N__39095\,
            I => \N__39026\
        );

    \I__9947\ : InMux
    port map (
            O => \N__39094\,
            I => \N__39023\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__39091\,
            I => \N__39020\
        );

    \I__9945\ : Span4Mux_s2_h
    port map (
            O => \N__39088\,
            I => \N__39015\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__39085\,
            I => \N__39015\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__39082\,
            I => \N__39012\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__39079\,
            I => \N__39007\
        );

    \I__9941\ : Span4Mux_h
    port map (
            O => \N__39074\,
            I => \N__39007\
        );

    \I__9940\ : Span4Mux_h
    port map (
            O => \N__39071\,
            I => \N__39000\
        );

    \I__9939\ : Span4Mux_v
    port map (
            O => \N__39068\,
            I => \N__39000\
        );

    \I__9938\ : Span4Mux_h
    port map (
            O => \N__39059\,
            I => \N__39000\
        );

    \I__9937\ : Span4Mux_h
    port map (
            O => \N__39056\,
            I => \N__38995\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__39053\,
            I => \N__38995\
        );

    \I__9935\ : InMux
    port map (
            O => \N__39052\,
            I => \N__38992\
        );

    \I__9934\ : Span12Mux_s6_h
    port map (
            O => \N__39049\,
            I => \N__38989\
        );

    \I__9933\ : Span4Mux_h
    port map (
            O => \N__39044\,
            I => \N__38982\
        );

    \I__9932\ : Span4Mux_h
    port map (
            O => \N__39039\,
            I => \N__38982\
        );

    \I__9931\ : Span4Mux_v
    port map (
            O => \N__39032\,
            I => \N__38982\
        );

    \I__9930\ : Span12Mux_s1_h
    port map (
            O => \N__39029\,
            I => \N__38977\
        );

    \I__9929\ : Span12Mux_s8_v
    port map (
            O => \N__39026\,
            I => \N__38977\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__39023\,
            I => \N__38970\
        );

    \I__9927\ : Span4Mux_h
    port map (
            O => \N__39020\,
            I => \N__38970\
        );

    \I__9926\ : Span4Mux_h
    port map (
            O => \N__39015\,
            I => \N__38970\
        );

    \I__9925\ : Span12Mux_s5_h
    port map (
            O => \N__39012\,
            I => \N__38961\
        );

    \I__9924\ : Sp12to4
    port map (
            O => \N__39007\,
            I => \N__38961\
        );

    \I__9923\ : Sp12to4
    port map (
            O => \N__39000\,
            I => \N__38961\
        );

    \I__9922\ : Sp12to4
    port map (
            O => \N__38995\,
            I => \N__38961\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__38992\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\
        );

    \I__9920\ : Odrv12
    port map (
            O => \N__38989\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\
        );

    \I__9919\ : Odrv4
    port map (
            O => \N__38982\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\
        );

    \I__9918\ : Odrv12
    port map (
            O => \N__38977\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__38970\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\
        );

    \I__9916\ : Odrv12
    port map (
            O => \N__38961\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\
        );

    \I__9915\ : CascadeMux
    port map (
            O => \N__38948\,
            I => \N__38945\
        );

    \I__9914\ : InMux
    port map (
            O => \N__38945\,
            I => \N__38942\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__38942\,
            I => \N__38938\
        );

    \I__9912\ : InMux
    port map (
            O => \N__38941\,
            I => \N__38935\
        );

    \I__9911\ : Span4Mux_v
    port map (
            O => \N__38938\,
            I => \N__38932\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__38935\,
            I => \N__38929\
        );

    \I__9909\ : Odrv4
    port map (
            O => \N__38932\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1\
        );

    \I__9908\ : Odrv12
    port map (
            O => \N__38929\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1\
        );

    \I__9907\ : InMux
    port map (
            O => \N__38924\,
            I => \N__38921\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__38921\,
            I => \N__38917\
        );

    \I__9905\ : InMux
    port map (
            O => \N__38920\,
            I => \N__38914\
        );

    \I__9904\ : Odrv4
    port map (
            O => \N__38917\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__38914\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1\
        );

    \I__9902\ : CascadeMux
    port map (
            O => \N__38909\,
            I => \N__38906\
        );

    \I__9901\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38903\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__38903\,
            I => \N__38900\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__38900\,
            I => \N__38897\
        );

    \I__9898\ : Span4Mux_s0_h
    port map (
            O => \N__38897\,
            I => \N__38894\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__38894\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_1\
        );

    \I__9896\ : CascadeMux
    port map (
            O => \N__38891\,
            I => \N__38883\
        );

    \I__9895\ : CascadeMux
    port map (
            O => \N__38890\,
            I => \N__38875\
        );

    \I__9894\ : InMux
    port map (
            O => \N__38889\,
            I => \N__38871\
        );

    \I__9893\ : CascadeMux
    port map (
            O => \N__38888\,
            I => \N__38868\
        );

    \I__9892\ : InMux
    port map (
            O => \N__38887\,
            I => \N__38864\
        );

    \I__9891\ : InMux
    port map (
            O => \N__38886\,
            I => \N__38861\
        );

    \I__9890\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38858\
        );

    \I__9889\ : InMux
    port map (
            O => \N__38882\,
            I => \N__38855\
        );

    \I__9888\ : CascadeMux
    port map (
            O => \N__38881\,
            I => \N__38852\
        );

    \I__9887\ : CascadeMux
    port map (
            O => \N__38880\,
            I => \N__38848\
        );

    \I__9886\ : CascadeMux
    port map (
            O => \N__38879\,
            I => \N__38844\
        );

    \I__9885\ : InMux
    port map (
            O => \N__38878\,
            I => \N__38840\
        );

    \I__9884\ : InMux
    port map (
            O => \N__38875\,
            I => \N__38837\
        );

    \I__9883\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38827\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__38871\,
            I => \N__38824\
        );

    \I__9881\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38821\
        );

    \I__9880\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38817\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__38864\,
            I => \N__38814\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__38861\,
            I => \N__38811\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__38858\,
            I => \N__38806\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__38855\,
            I => \N__38806\
        );

    \I__9875\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38803\
        );

    \I__9874\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38796\
        );

    \I__9873\ : InMux
    port map (
            O => \N__38848\,
            I => \N__38793\
        );

    \I__9872\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38790\
        );

    \I__9871\ : InMux
    port map (
            O => \N__38844\,
            I => \N__38787\
        );

    \I__9870\ : CascadeMux
    port map (
            O => \N__38843\,
            I => \N__38784\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__38840\,
            I => \N__38779\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__38837\,
            I => \N__38776\
        );

    \I__9867\ : InMux
    port map (
            O => \N__38836\,
            I => \N__38773\
        );

    \I__9866\ : InMux
    port map (
            O => \N__38835\,
            I => \N__38770\
        );

    \I__9865\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38767\
        );

    \I__9864\ : CascadeMux
    port map (
            O => \N__38833\,
            I => \N__38764\
        );

    \I__9863\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38761\
        );

    \I__9862\ : InMux
    port map (
            O => \N__38831\,
            I => \N__38758\
        );

    \I__9861\ : InMux
    port map (
            O => \N__38830\,
            I => \N__38755\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__38827\,
            I => \N__38752\
        );

    \I__9859\ : Span4Mux_v
    port map (
            O => \N__38824\,
            I => \N__38747\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__38821\,
            I => \N__38747\
        );

    \I__9857\ : InMux
    port map (
            O => \N__38820\,
            I => \N__38744\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__38817\,
            I => \N__38739\
        );

    \I__9855\ : Span4Mux_s3_h
    port map (
            O => \N__38814\,
            I => \N__38739\
        );

    \I__9854\ : Span4Mux_v
    port map (
            O => \N__38811\,
            I => \N__38732\
        );

    \I__9853\ : Span4Mux_s3_h
    port map (
            O => \N__38806\,
            I => \N__38732\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__38803\,
            I => \N__38732\
        );

    \I__9851\ : CascadeMux
    port map (
            O => \N__38802\,
            I => \N__38726\
        );

    \I__9850\ : InMux
    port map (
            O => \N__38801\,
            I => \N__38722\
        );

    \I__9849\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38719\
        );

    \I__9848\ : InMux
    port map (
            O => \N__38799\,
            I => \N__38716\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__38796\,
            I => \N__38711\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__38793\,
            I => \N__38711\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__38790\,
            I => \N__38706\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__38787\,
            I => \N__38706\
        );

    \I__9843\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38703\
        );

    \I__9842\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38700\
        );

    \I__9841\ : InMux
    port map (
            O => \N__38782\,
            I => \N__38697\
        );

    \I__9840\ : Span4Mux_h
    port map (
            O => \N__38779\,
            I => \N__38686\
        );

    \I__9839\ : Span4Mux_s3_h
    port map (
            O => \N__38776\,
            I => \N__38686\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__38773\,
            I => \N__38686\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__38770\,
            I => \N__38686\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__38767\,
            I => \N__38686\
        );

    \I__9835\ : InMux
    port map (
            O => \N__38764\,
            I => \N__38683\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__38761\,
            I => \N__38678\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__38758\,
            I => \N__38678\
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__38755\,
            I => \N__38673\
        );

    \I__9831\ : Span4Mux_s2_v
    port map (
            O => \N__38752\,
            I => \N__38673\
        );

    \I__9830\ : Span4Mux_s1_h
    port map (
            O => \N__38747\,
            I => \N__38670\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__38744\,
            I => \N__38663\
        );

    \I__9828\ : Span4Mux_v
    port map (
            O => \N__38739\,
            I => \N__38663\
        );

    \I__9827\ : Span4Mux_h
    port map (
            O => \N__38732\,
            I => \N__38663\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__38731\,
            I => \N__38660\
        );

    \I__9825\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38657\
        );

    \I__9824\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38654\
        );

    \I__9823\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38651\
        );

    \I__9822\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38648\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__38722\,
            I => \N__38641\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__38719\,
            I => \N__38641\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__38716\,
            I => \N__38641\
        );

    \I__9818\ : Span4Mux_v
    port map (
            O => \N__38711\,
            I => \N__38636\
        );

    \I__9817\ : Span4Mux_s2_v
    port map (
            O => \N__38706\,
            I => \N__38636\
        );

    \I__9816\ : LocalMux
    port map (
            O => \N__38703\,
            I => \N__38633\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__38700\,
            I => \N__38626\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__38697\,
            I => \N__38626\
        );

    \I__9813\ : Sp12to4
    port map (
            O => \N__38686\,
            I => \N__38626\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__38683\,
            I => \N__38617\
        );

    \I__9811\ : Span4Mux_v
    port map (
            O => \N__38678\,
            I => \N__38617\
        );

    \I__9810\ : Span4Mux_v
    port map (
            O => \N__38673\,
            I => \N__38617\
        );

    \I__9809\ : Span4Mux_v
    port map (
            O => \N__38670\,
            I => \N__38617\
        );

    \I__9808\ : Sp12to4
    port map (
            O => \N__38663\,
            I => \N__38614\
        );

    \I__9807\ : InMux
    port map (
            O => \N__38660\,
            I => \N__38611\
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__38657\,
            I => \N__38604\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38604\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__38651\,
            I => \N__38604\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__38648\,
            I => \N__38599\
        );

    \I__9802\ : Span12Mux_s10_h
    port map (
            O => \N__38641\,
            I => \N__38599\
        );

    \I__9801\ : Span4Mux_v
    port map (
            O => \N__38636\,
            I => \N__38596\
        );

    \I__9800\ : Span12Mux_s3_h
    port map (
            O => \N__38633\,
            I => \N__38585\
        );

    \I__9799\ : Span12Mux_s6_v
    port map (
            O => \N__38626\,
            I => \N__38585\
        );

    \I__9798\ : Sp12to4
    port map (
            O => \N__38617\,
            I => \N__38585\
        );

    \I__9797\ : Span12Mux_s9_v
    port map (
            O => \N__38614\,
            I => \N__38585\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__38611\,
            I => \N__38585\
        );

    \I__9795\ : Odrv12
    port map (
            O => \N__38604\,
            I => \processor_zipi8.arith_logical_result_2\
        );

    \I__9794\ : Odrv12
    port map (
            O => \N__38599\,
            I => \processor_zipi8.arith_logical_result_2\
        );

    \I__9793\ : Odrv4
    port map (
            O => \N__38596\,
            I => \processor_zipi8.arith_logical_result_2\
        );

    \I__9792\ : Odrv12
    port map (
            O => \N__38585\,
            I => \processor_zipi8.arith_logical_result_2\
        );

    \I__9791\ : CascadeMux
    port map (
            O => \N__38576\,
            I => \N__38571\
        );

    \I__9790\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38562\
        );

    \I__9789\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38559\
        );

    \I__9788\ : InMux
    port map (
            O => \N__38571\,
            I => \N__38553\
        );

    \I__9787\ : CascadeMux
    port map (
            O => \N__38570\,
            I => \N__38546\
        );

    \I__9786\ : CascadeMux
    port map (
            O => \N__38569\,
            I => \N__38542\
        );

    \I__9785\ : CascadeMux
    port map (
            O => \N__38568\,
            I => \N__38537\
        );

    \I__9784\ : CascadeMux
    port map (
            O => \N__38567\,
            I => \N__38534\
        );

    \I__9783\ : InMux
    port map (
            O => \N__38566\,
            I => \N__38527\
        );

    \I__9782\ : InMux
    port map (
            O => \N__38565\,
            I => \N__38524\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__38562\,
            I => \N__38519\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__38559\,
            I => \N__38519\
        );

    \I__9779\ : CascadeMux
    port map (
            O => \N__38558\,
            I => \N__38514\
        );

    \I__9778\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38510\
        );

    \I__9777\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38507\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__38553\,
            I => \N__38502\
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__38552\,
            I => \N__38499\
        );

    \I__9774\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38496\
        );

    \I__9773\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38493\
        );

    \I__9772\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38490\
        );

    \I__9771\ : InMux
    port map (
            O => \N__38546\,
            I => \N__38487\
        );

    \I__9770\ : InMux
    port map (
            O => \N__38545\,
            I => \N__38484\
        );

    \I__9769\ : InMux
    port map (
            O => \N__38542\,
            I => \N__38481\
        );

    \I__9768\ : InMux
    port map (
            O => \N__38541\,
            I => \N__38478\
        );

    \I__9767\ : CascadeMux
    port map (
            O => \N__38540\,
            I => \N__38475\
        );

    \I__9766\ : InMux
    port map (
            O => \N__38537\,
            I => \N__38472\
        );

    \I__9765\ : InMux
    port map (
            O => \N__38534\,
            I => \N__38469\
        );

    \I__9764\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38466\
        );

    \I__9763\ : CascadeMux
    port map (
            O => \N__38532\,
            I => \N__38463\
        );

    \I__9762\ : CascadeMux
    port map (
            O => \N__38531\,
            I => \N__38458\
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__38530\,
            I => \N__38455\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__38527\,
            I => \N__38452\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__38524\,
            I => \N__38447\
        );

    \I__9758\ : Span4Mux_v
    port map (
            O => \N__38519\,
            I => \N__38447\
        );

    \I__9757\ : CascadeMux
    port map (
            O => \N__38518\,
            I => \N__38443\
        );

    \I__9756\ : CascadeMux
    port map (
            O => \N__38517\,
            I => \N__38440\
        );

    \I__9755\ : InMux
    port map (
            O => \N__38514\,
            I => \N__38437\
        );

    \I__9754\ : InMux
    port map (
            O => \N__38513\,
            I => \N__38434\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__38510\,
            I => \N__38429\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__38507\,
            I => \N__38429\
        );

    \I__9751\ : CascadeMux
    port map (
            O => \N__38506\,
            I => \N__38426\
        );

    \I__9750\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38422\
        );

    \I__9749\ : Span4Mux_v
    port map (
            O => \N__38502\,
            I => \N__38419\
        );

    \I__9748\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38416\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__38496\,
            I => \N__38411\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__38493\,
            I => \N__38411\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__38490\,
            I => \N__38406\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__38487\,
            I => \N__38406\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__38484\,
            I => \N__38403\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__38481\,
            I => \N__38398\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__38478\,
            I => \N__38398\
        );

    \I__9740\ : InMux
    port map (
            O => \N__38475\,
            I => \N__38395\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__38472\,
            I => \N__38388\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__38469\,
            I => \N__38388\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__38466\,
            I => \N__38388\
        );

    \I__9736\ : InMux
    port map (
            O => \N__38463\,
            I => \N__38385\
        );

    \I__9735\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38382\
        );

    \I__9734\ : CascadeMux
    port map (
            O => \N__38461\,
            I => \N__38379\
        );

    \I__9733\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38376\
        );

    \I__9732\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38373\
        );

    \I__9731\ : Span4Mux_v
    port map (
            O => \N__38452\,
            I => \N__38368\
        );

    \I__9730\ : Span4Mux_v
    port map (
            O => \N__38447\,
            I => \N__38368\
        );

    \I__9729\ : InMux
    port map (
            O => \N__38446\,
            I => \N__38365\
        );

    \I__9728\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38362\
        );

    \I__9727\ : InMux
    port map (
            O => \N__38440\,
            I => \N__38359\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__38437\,
            I => \N__38352\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__38434\,
            I => \N__38352\
        );

    \I__9724\ : Span4Mux_v
    port map (
            O => \N__38429\,
            I => \N__38352\
        );

    \I__9723\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38349\
        );

    \I__9722\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38346\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__38422\,
            I => \N__38341\
        );

    \I__9720\ : Span4Mux_v
    port map (
            O => \N__38419\,
            I => \N__38341\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38334\
        );

    \I__9718\ : Span4Mux_v
    port map (
            O => \N__38411\,
            I => \N__38334\
        );

    \I__9717\ : Span4Mux_s3_h
    port map (
            O => \N__38406\,
            I => \N__38334\
        );

    \I__9716\ : Span4Mux_v
    port map (
            O => \N__38403\,
            I => \N__38325\
        );

    \I__9715\ : Span4Mux_s3_h
    port map (
            O => \N__38398\,
            I => \N__38325\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__38395\,
            I => \N__38325\
        );

    \I__9713\ : Span4Mux_v
    port map (
            O => \N__38388\,
            I => \N__38325\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__38385\,
            I => \N__38320\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__38382\,
            I => \N__38320\
        );

    \I__9710\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38317\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__38376\,
            I => \N__38314\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__38373\,
            I => \N__38311\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__38368\,
            I => \N__38307\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__38365\,
            I => \N__38302\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__38362\,
            I => \N__38302\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__38359\,
            I => \N__38299\
        );

    \I__9703\ : Span4Mux_v
    port map (
            O => \N__38352\,
            I => \N__38296\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__38349\,
            I => \N__38289\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__38346\,
            I => \N__38289\
        );

    \I__9700\ : Span4Mux_v
    port map (
            O => \N__38341\,
            I => \N__38289\
        );

    \I__9699\ : Span4Mux_h
    port map (
            O => \N__38334\,
            I => \N__38282\
        );

    \I__9698\ : Span4Mux_h
    port map (
            O => \N__38325\,
            I => \N__38282\
        );

    \I__9697\ : Span4Mux_v
    port map (
            O => \N__38320\,
            I => \N__38282\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__38317\,
            I => \N__38279\
        );

    \I__9695\ : Span4Mux_s3_v
    port map (
            O => \N__38314\,
            I => \N__38274\
        );

    \I__9694\ : Span4Mux_v
    port map (
            O => \N__38311\,
            I => \N__38274\
        );

    \I__9693\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38271\
        );

    \I__9692\ : Span4Mux_h
    port map (
            O => \N__38307\,
            I => \N__38268\
        );

    \I__9691\ : Span4Mux_s2_v
    port map (
            O => \N__38302\,
            I => \N__38259\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__38299\,
            I => \N__38259\
        );

    \I__9689\ : Span4Mux_v
    port map (
            O => \N__38296\,
            I => \N__38259\
        );

    \I__9688\ : Span4Mux_h
    port map (
            O => \N__38289\,
            I => \N__38259\
        );

    \I__9687\ : Span4Mux_v
    port map (
            O => \N__38282\,
            I => \N__38256\
        );

    \I__9686\ : Span4Mux_h
    port map (
            O => \N__38279\,
            I => \N__38249\
        );

    \I__9685\ : Span4Mux_h
    port map (
            O => \N__38274\,
            I => \N__38249\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__38271\,
            I => \N__38249\
        );

    \I__9683\ : Odrv4
    port map (
            O => \N__38268\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265\
        );

    \I__9682\ : Odrv4
    port map (
            O => \N__38259\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265\
        );

    \I__9681\ : Odrv4
    port map (
            O => \N__38256\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265\
        );

    \I__9680\ : Odrv4
    port map (
            O => \N__38249\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265\
        );

    \I__9679\ : InMux
    port map (
            O => \N__38240\,
            I => \N__38237\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__38237\,
            I => \N__38233\
        );

    \I__9677\ : InMux
    port map (
            O => \N__38236\,
            I => \N__38230\
        );

    \I__9676\ : Span4Mux_s3_h
    port map (
            O => \N__38233\,
            I => \N__38227\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__38230\,
            I => \N__38224\
        );

    \I__9674\ : Odrv4
    port map (
            O => \N__38227\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2\
        );

    \I__9673\ : Odrv12
    port map (
            O => \N__38224\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2\
        );

    \I__9672\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38216\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__38216\,
            I => \N__38212\
        );

    \I__9670\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38209\
        );

    \I__9669\ : Odrv4
    port map (
            O => \N__38212\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__38209\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2\
        );

    \I__9667\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38201\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__38201\,
            I => \N__38198\
        );

    \I__9665\ : Span4Mux_h
    port map (
            O => \N__38198\,
            I => \N__38195\
        );

    \I__9664\ : Odrv4
    port map (
            O => \N__38195\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_2\
        );

    \I__9663\ : CascadeMux
    port map (
            O => \N__38192\,
            I => \N__38178\
        );

    \I__9662\ : CascadeMux
    port map (
            O => \N__38191\,
            I => \N__38175\
        );

    \I__9661\ : CascadeMux
    port map (
            O => \N__38190\,
            I => \N__38169\
        );

    \I__9660\ : CascadeMux
    port map (
            O => \N__38189\,
            I => \N__38166\
        );

    \I__9659\ : CascadeMux
    port map (
            O => \N__38188\,
            I => \N__38163\
        );

    \I__9658\ : CascadeMux
    port map (
            O => \N__38187\,
            I => \N__38160\
        );

    \I__9657\ : CascadeMux
    port map (
            O => \N__38186\,
            I => \N__38155\
        );

    \I__9656\ : CascadeMux
    port map (
            O => \N__38185\,
            I => \N__38151\
        );

    \I__9655\ : CascadeMux
    port map (
            O => \N__38184\,
            I => \N__38148\
        );

    \I__9654\ : CascadeMux
    port map (
            O => \N__38183\,
            I => \N__38141\
        );

    \I__9653\ : CascadeMux
    port map (
            O => \N__38182\,
            I => \N__38138\
        );

    \I__9652\ : CascadeMux
    port map (
            O => \N__38181\,
            I => \N__38133\
        );

    \I__9651\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38130\
        );

    \I__9650\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38127\
        );

    \I__9649\ : CascadeMux
    port map (
            O => \N__38174\,
            I => \N__38124\
        );

    \I__9648\ : CascadeMux
    port map (
            O => \N__38173\,
            I => \N__38119\
        );

    \I__9647\ : CascadeMux
    port map (
            O => \N__38172\,
            I => \N__38115\
        );

    \I__9646\ : InMux
    port map (
            O => \N__38169\,
            I => \N__38112\
        );

    \I__9645\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38109\
        );

    \I__9644\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38106\
        );

    \I__9643\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38103\
        );

    \I__9642\ : CascadeMux
    port map (
            O => \N__38159\,
            I => \N__38100\
        );

    \I__9641\ : CascadeMux
    port map (
            O => \N__38158\,
            I => \N__38095\
        );

    \I__9640\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38092\
        );

    \I__9639\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38089\
        );

    \I__9638\ : InMux
    port map (
            O => \N__38151\,
            I => \N__38086\
        );

    \I__9637\ : InMux
    port map (
            O => \N__38148\,
            I => \N__38083\
        );

    \I__9636\ : InMux
    port map (
            O => \N__38147\,
            I => \N__38080\
        );

    \I__9635\ : CascadeMux
    port map (
            O => \N__38146\,
            I => \N__38075\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__38145\,
            I => \N__38072\
        );

    \I__9633\ : InMux
    port map (
            O => \N__38144\,
            I => \N__38068\
        );

    \I__9632\ : InMux
    port map (
            O => \N__38141\,
            I => \N__38064\
        );

    \I__9631\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38061\
        );

    \I__9630\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38058\
        );

    \I__9629\ : InMux
    port map (
            O => \N__38136\,
            I => \N__38055\
        );

    \I__9628\ : InMux
    port map (
            O => \N__38133\,
            I => \N__38052\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__38130\,
            I => \N__38047\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__38127\,
            I => \N__38047\
        );

    \I__9625\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38044\
        );

    \I__9624\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38041\
        );

    \I__9623\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38038\
        );

    \I__9622\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38035\
        );

    \I__9621\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38032\
        );

    \I__9620\ : InMux
    port map (
            O => \N__38115\,
            I => \N__38029\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__38112\,
            I => \N__38026\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__38109\,
            I => \N__38019\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__38106\,
            I => \N__38019\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__38103\,
            I => \N__38019\
        );

    \I__9615\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38016\
        );

    \I__9614\ : InMux
    port map (
            O => \N__38099\,
            I => \N__38013\
        );

    \I__9613\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38010\
        );

    \I__9612\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38007\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__38092\,
            I => \N__38004\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__38089\,
            I => \N__37995\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__38086\,
            I => \N__37995\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__38083\,
            I => \N__37995\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__37995\
        );

    \I__9606\ : InMux
    port map (
            O => \N__38079\,
            I => \N__37992\
        );

    \I__9605\ : InMux
    port map (
            O => \N__38078\,
            I => \N__37989\
        );

    \I__9604\ : InMux
    port map (
            O => \N__38075\,
            I => \N__37986\
        );

    \I__9603\ : InMux
    port map (
            O => \N__38072\,
            I => \N__37983\
        );

    \I__9602\ : InMux
    port map (
            O => \N__38071\,
            I => \N__37980\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__38068\,
            I => \N__37977\
        );

    \I__9600\ : InMux
    port map (
            O => \N__38067\,
            I => \N__37974\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__38064\,
            I => \N__37969\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__38061\,
            I => \N__37969\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__38058\,
            I => \N__37960\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__38055\,
            I => \N__37960\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__38052\,
            I => \N__37960\
        );

    \I__9594\ : Span4Mux_v
    port map (
            O => \N__38047\,
            I => \N__37960\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__38044\,
            I => \N__37957\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__38041\,
            I => \N__37954\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__38038\,
            I => \N__37951\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__38035\,
            I => \N__37948\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__38032\,
            I => \N__37939\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__38029\,
            I => \N__37939\
        );

    \I__9587\ : Span4Mux_s3_h
    port map (
            O => \N__38026\,
            I => \N__37939\
        );

    \I__9586\ : Span4Mux_v
    port map (
            O => \N__38019\,
            I => \N__37939\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__38016\,
            I => \N__37936\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__38013\,
            I => \N__37929\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__38010\,
            I => \N__37929\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__38007\,
            I => \N__37929\
        );

    \I__9581\ : Span4Mux_v
    port map (
            O => \N__38004\,
            I => \N__37926\
        );

    \I__9580\ : Span4Mux_v
    port map (
            O => \N__37995\,
            I => \N__37923\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__37992\,
            I => \N__37910\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__37989\,
            I => \N__37910\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37910\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37910\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__37980\,
            I => \N__37910\
        );

    \I__9574\ : Span4Mux_s2_v
    port map (
            O => \N__37977\,
            I => \N__37910\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__37974\,
            I => \N__37903\
        );

    \I__9572\ : Span4Mux_v
    port map (
            O => \N__37969\,
            I => \N__37903\
        );

    \I__9571\ : Span4Mux_v
    port map (
            O => \N__37960\,
            I => \N__37903\
        );

    \I__9570\ : Span4Mux_s3_h
    port map (
            O => \N__37957\,
            I => \N__37900\
        );

    \I__9569\ : Span4Mux_v
    port map (
            O => \N__37954\,
            I => \N__37890\
        );

    \I__9568\ : Span4Mux_s3_h
    port map (
            O => \N__37951\,
            I => \N__37890\
        );

    \I__9567\ : Span4Mux_v
    port map (
            O => \N__37948\,
            I => \N__37890\
        );

    \I__9566\ : Span4Mux_v
    port map (
            O => \N__37939\,
            I => \N__37890\
        );

    \I__9565\ : Span4Mux_v
    port map (
            O => \N__37936\,
            I => \N__37881\
        );

    \I__9564\ : Span4Mux_v
    port map (
            O => \N__37929\,
            I => \N__37881\
        );

    \I__9563\ : Span4Mux_h
    port map (
            O => \N__37926\,
            I => \N__37881\
        );

    \I__9562\ : Span4Mux_h
    port map (
            O => \N__37923\,
            I => \N__37881\
        );

    \I__9561\ : Span4Mux_v
    port map (
            O => \N__37910\,
            I => \N__37874\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__37903\,
            I => \N__37874\
        );

    \I__9559\ : Span4Mux_v
    port map (
            O => \N__37900\,
            I => \N__37874\
        );

    \I__9558\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37871\
        );

    \I__9557\ : Odrv4
    port map (
            O => \N__37890\,
            I => \processor_zipi8.arith_logical_result_3\
        );

    \I__9556\ : Odrv4
    port map (
            O => \N__37881\,
            I => \processor_zipi8.arith_logical_result_3\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__37874\,
            I => \processor_zipi8.arith_logical_result_3\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__37871\,
            I => \processor_zipi8.arith_logical_result_3\
        );

    \I__9553\ : CascadeMux
    port map (
            O => \N__37862\,
            I => \N__37859\
        );

    \I__9552\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37854\
        );

    \I__9551\ : CascadeMux
    port map (
            O => \N__37858\,
            I => \N__37850\
        );

    \I__9550\ : CascadeMux
    port map (
            O => \N__37857\,
            I => \N__37847\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__37854\,
            I => \N__37844\
        );

    \I__9548\ : CascadeMux
    port map (
            O => \N__37853\,
            I => \N__37841\
        );

    \I__9547\ : InMux
    port map (
            O => \N__37850\,
            I => \N__37837\
        );

    \I__9546\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37832\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__37844\,
            I => \N__37829\
        );

    \I__9544\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37826\
        );

    \I__9543\ : CascadeMux
    port map (
            O => \N__37840\,
            I => \N__37820\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__37837\,
            I => \N__37817\
        );

    \I__9541\ : InMux
    port map (
            O => \N__37836\,
            I => \N__37814\
        );

    \I__9540\ : CascadeMux
    port map (
            O => \N__37835\,
            I => \N__37811\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__37832\,
            I => \N__37807\
        );

    \I__9538\ : Span4Mux_h
    port map (
            O => \N__37829\,
            I => \N__37802\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__37826\,
            I => \N__37802\
        );

    \I__9536\ : InMux
    port map (
            O => \N__37825\,
            I => \N__37798\
        );

    \I__9535\ : CascadeMux
    port map (
            O => \N__37824\,
            I => \N__37794\
        );

    \I__9534\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37790\
        );

    \I__9533\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37787\
        );

    \I__9532\ : Span4Mux_s0_h
    port map (
            O => \N__37817\,
            I => \N__37782\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37782\
        );

    \I__9530\ : InMux
    port map (
            O => \N__37811\,
            I => \N__37779\
        );

    \I__9529\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37775\
        );

    \I__9528\ : Span4Mux_h
    port map (
            O => \N__37807\,
            I => \N__37769\
        );

    \I__9527\ : Span4Mux_v
    port map (
            O => \N__37802\,
            I => \N__37769\
        );

    \I__9526\ : InMux
    port map (
            O => \N__37801\,
            I => \N__37766\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__37798\,
            I => \N__37763\
        );

    \I__9524\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37760\
        );

    \I__9523\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37757\
        );

    \I__9522\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37750\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__37790\,
            I => \N__37741\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__37787\,
            I => \N__37741\
        );

    \I__9519\ : Span4Mux_v
    port map (
            O => \N__37782\,
            I => \N__37741\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__37779\,
            I => \N__37741\
        );

    \I__9517\ : InMux
    port map (
            O => \N__37778\,
            I => \N__37738\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__37775\,
            I => \N__37735\
        );

    \I__9515\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37732\
        );

    \I__9514\ : Span4Mux_v
    port map (
            O => \N__37769\,
            I => \N__37727\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__37766\,
            I => \N__37727\
        );

    \I__9512\ : Span4Mux_v
    port map (
            O => \N__37763\,
            I => \N__37722\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__37760\,
            I => \N__37722\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37719\
        );

    \I__9509\ : InMux
    port map (
            O => \N__37756\,
            I => \N__37716\
        );

    \I__9508\ : InMux
    port map (
            O => \N__37755\,
            I => \N__37713\
        );

    \I__9507\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37710\
        );

    \I__9506\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37707\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37698\
        );

    \I__9504\ : Span4Mux_v
    port map (
            O => \N__37741\,
            I => \N__37693\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__37738\,
            I => \N__37693\
        );

    \I__9502\ : Span4Mux_v
    port map (
            O => \N__37735\,
            I => \N__37690\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__37732\,
            I => \N__37685\
        );

    \I__9500\ : Span4Mux_v
    port map (
            O => \N__37727\,
            I => \N__37685\
        );

    \I__9499\ : Span4Mux_v
    port map (
            O => \N__37722\,
            I => \N__37680\
        );

    \I__9498\ : Span4Mux_v
    port map (
            O => \N__37719\,
            I => \N__37680\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37677\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__37713\,
            I => \N__37674\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__37710\,
            I => \N__37669\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__37707\,
            I => \N__37669\
        );

    \I__9493\ : CascadeMux
    port map (
            O => \N__37706\,
            I => \N__37665\
        );

    \I__9492\ : InMux
    port map (
            O => \N__37705\,
            I => \N__37662\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__37704\,
            I => \N__37658\
        );

    \I__9490\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37655\
        );

    \I__9489\ : InMux
    port map (
            O => \N__37702\,
            I => \N__37651\
        );

    \I__9488\ : InMux
    port map (
            O => \N__37701\,
            I => \N__37648\
        );

    \I__9487\ : Span4Mux_v
    port map (
            O => \N__37698\,
            I => \N__37641\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__37693\,
            I => \N__37641\
        );

    \I__9485\ : Span4Mux_s0_h
    port map (
            O => \N__37690\,
            I => \N__37641\
        );

    \I__9484\ : Span4Mux_h
    port map (
            O => \N__37685\,
            I => \N__37630\
        );

    \I__9483\ : Span4Mux_h
    port map (
            O => \N__37680\,
            I => \N__37630\
        );

    \I__9482\ : Span4Mux_s2_h
    port map (
            O => \N__37677\,
            I => \N__37630\
        );

    \I__9481\ : Span4Mux_v
    port map (
            O => \N__37674\,
            I => \N__37630\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__37669\,
            I => \N__37630\
        );

    \I__9479\ : CascadeMux
    port map (
            O => \N__37668\,
            I => \N__37624\
        );

    \I__9478\ : InMux
    port map (
            O => \N__37665\,
            I => \N__37621\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__37662\,
            I => \N__37618\
        );

    \I__9476\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37615\
        );

    \I__9475\ : InMux
    port map (
            O => \N__37658\,
            I => \N__37612\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__37655\,
            I => \N__37609\
        );

    \I__9473\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37606\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__37651\,
            I => \N__37603\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__37648\,
            I => \N__37600\
        );

    \I__9470\ : Sp12to4
    port map (
            O => \N__37641\,
            I => \N__37595\
        );

    \I__9469\ : Sp12to4
    port map (
            O => \N__37630\,
            I => \N__37595\
        );

    \I__9468\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37592\
        );

    \I__9467\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37589\
        );

    \I__9466\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37586\
        );

    \I__9465\ : InMux
    port map (
            O => \N__37624\,
            I => \N__37583\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__37621\,
            I => \N__37580\
        );

    \I__9463\ : Span4Mux_s2_v
    port map (
            O => \N__37618\,
            I => \N__37577\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__37615\,
            I => \N__37570\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__37612\,
            I => \N__37570\
        );

    \I__9460\ : Span4Mux_v
    port map (
            O => \N__37609\,
            I => \N__37570\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__37606\,
            I => \N__37565\
        );

    \I__9458\ : Span4Mux_v
    port map (
            O => \N__37603\,
            I => \N__37565\
        );

    \I__9457\ : Span12Mux_s6_h
    port map (
            O => \N__37600\,
            I => \N__37560\
        );

    \I__9456\ : Span12Mux_s5_h
    port map (
            O => \N__37595\,
            I => \N__37560\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__37592\,
            I => \N__37555\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__37589\,
            I => \N__37555\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__37586\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__37583\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__37580\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9450\ : Odrv4
    port map (
            O => \N__37577\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9449\ : Odrv4
    port map (
            O => \N__37570\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9448\ : Odrv4
    port map (
            O => \N__37565\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9447\ : Odrv12
    port map (
            O => \N__37560\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9446\ : Odrv12
    port map (
            O => \N__37555\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\
        );

    \I__9445\ : InMux
    port map (
            O => \N__37538\,
            I => \N__37535\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__37535\,
            I => \N__37531\
        );

    \I__9443\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37528\
        );

    \I__9442\ : Span4Mux_v
    port map (
            O => \N__37531\,
            I => \N__37523\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__37528\,
            I => \N__37523\
        );

    \I__9440\ : Span4Mux_s0_h
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__9439\ : Odrv4
    port map (
            O => \N__37520\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_3\
        );

    \I__9438\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37513\
        );

    \I__9437\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37510\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__37513\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__37510\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3\
        );

    \I__9434\ : InMux
    port map (
            O => \N__37505\,
            I => \N__37491\
        );

    \I__9433\ : InMux
    port map (
            O => \N__37504\,
            I => \N__37479\
        );

    \I__9432\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37479\
        );

    \I__9431\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37470\
        );

    \I__9430\ : InMux
    port map (
            O => \N__37501\,
            I => \N__37470\
        );

    \I__9429\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37470\
        );

    \I__9428\ : InMux
    port map (
            O => \N__37499\,
            I => \N__37462\
        );

    \I__9427\ : InMux
    port map (
            O => \N__37498\,
            I => \N__37462\
        );

    \I__9426\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37457\
        );

    \I__9425\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37457\
        );

    \I__9424\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37452\
        );

    \I__9423\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37452\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__37491\,
            I => \N__37445\
        );

    \I__9421\ : InMux
    port map (
            O => \N__37490\,
            I => \N__37442\
        );

    \I__9420\ : InMux
    port map (
            O => \N__37489\,
            I => \N__37433\
        );

    \I__9419\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37433\
        );

    \I__9418\ : InMux
    port map (
            O => \N__37487\,
            I => \N__37420\
        );

    \I__9417\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37417\
        );

    \I__9416\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37412\
        );

    \I__9415\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37412\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__37479\,
            I => \N__37406\
        );

    \I__9413\ : InMux
    port map (
            O => \N__37478\,
            I => \N__37401\
        );

    \I__9412\ : InMux
    port map (
            O => \N__37477\,
            I => \N__37401\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__37470\,
            I => \N__37398\
        );

    \I__9410\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37391\
        );

    \I__9409\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37386\
        );

    \I__9408\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37386\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__37462\,
            I => \N__37378\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__37457\,
            I => \N__37373\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__37452\,
            I => \N__37373\
        );

    \I__9404\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37369\
        );

    \I__9403\ : InMux
    port map (
            O => \N__37450\,
            I => \N__37362\
        );

    \I__9402\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37362\
        );

    \I__9401\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37362\
        );

    \I__9400\ : Span4Mux_v
    port map (
            O => \N__37445\,
            I => \N__37357\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__37442\,
            I => \N__37357\
        );

    \I__9398\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37349\
        );

    \I__9397\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37349\
        );

    \I__9396\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37346\
        );

    \I__9395\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37343\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__37433\,
            I => \N__37340\
        );

    \I__9393\ : InMux
    port map (
            O => \N__37432\,
            I => \N__37333\
        );

    \I__9392\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37333\
        );

    \I__9391\ : InMux
    port map (
            O => \N__37430\,
            I => \N__37333\
        );

    \I__9390\ : InMux
    port map (
            O => \N__37429\,
            I => \N__37324\
        );

    \I__9389\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37317\
        );

    \I__9388\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37317\
        );

    \I__9387\ : InMux
    port map (
            O => \N__37426\,
            I => \N__37310\
        );

    \I__9386\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37310\
        );

    \I__9385\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37310\
        );

    \I__9384\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37307\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__37420\,
            I => \N__37304\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__37417\,
            I => \N__37290\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__37412\,
            I => \N__37287\
        );

    \I__9380\ : InMux
    port map (
            O => \N__37411\,
            I => \N__37281\
        );

    \I__9379\ : InMux
    port map (
            O => \N__37410\,
            I => \N__37281\
        );

    \I__9378\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37278\
        );

    \I__9377\ : Span4Mux_s2_v
    port map (
            O => \N__37406\,
            I => \N__37273\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__37401\,
            I => \N__37273\
        );

    \I__9375\ : Span4Mux_v
    port map (
            O => \N__37398\,
            I => \N__37270\
        );

    \I__9374\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37265\
        );

    \I__9373\ : InMux
    port map (
            O => \N__37396\,
            I => \N__37265\
        );

    \I__9372\ : InMux
    port map (
            O => \N__37395\,
            I => \N__37260\
        );

    \I__9371\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37260\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__37391\,
            I => \N__37255\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__37386\,
            I => \N__37255\
        );

    \I__9368\ : CascadeMux
    port map (
            O => \N__37385\,
            I => \N__37246\
        );

    \I__9367\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37236\
        );

    \I__9366\ : InMux
    port map (
            O => \N__37383\,
            I => \N__37236\
        );

    \I__9365\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37236\
        );

    \I__9364\ : InMux
    port map (
            O => \N__37381\,
            I => \N__37236\
        );

    \I__9363\ : Span4Mux_v
    port map (
            O => \N__37378\,
            I => \N__37231\
        );

    \I__9362\ : Span4Mux_v
    port map (
            O => \N__37373\,
            I => \N__37231\
        );

    \I__9361\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37228\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__37369\,
            I => \N__37221\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__37362\,
            I => \N__37221\
        );

    \I__9358\ : Span4Mux_s3_v
    port map (
            O => \N__37357\,
            I => \N__37221\
        );

    \I__9357\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37218\
        );

    \I__9356\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37206\
        );

    \I__9355\ : InMux
    port map (
            O => \N__37354\,
            I => \N__37206\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__37349\,
            I => \N__37203\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__37346\,
            I => \N__37194\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__37343\,
            I => \N__37194\
        );

    \I__9351\ : Span4Mux_h
    port map (
            O => \N__37340\,
            I => \N__37194\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__37333\,
            I => \N__37194\
        );

    \I__9349\ : InMux
    port map (
            O => \N__37332\,
            I => \N__37183\
        );

    \I__9348\ : InMux
    port map (
            O => \N__37331\,
            I => \N__37183\
        );

    \I__9347\ : InMux
    port map (
            O => \N__37330\,
            I => \N__37183\
        );

    \I__9346\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37183\
        );

    \I__9345\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37183\
        );

    \I__9344\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37180\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__37324\,
            I => \N__37177\
        );

    \I__9342\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37172\
        );

    \I__9341\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37172\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37163\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__37310\,
            I => \N__37163\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__37307\,
            I => \N__37163\
        );

    \I__9337\ : Span4Mux_s3_v
    port map (
            O => \N__37304\,
            I => \N__37163\
        );

    \I__9336\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37154\
        );

    \I__9335\ : InMux
    port map (
            O => \N__37302\,
            I => \N__37154\
        );

    \I__9334\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37154\
        );

    \I__9333\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37154\
        );

    \I__9332\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37147\
        );

    \I__9331\ : InMux
    port map (
            O => \N__37298\,
            I => \N__37147\
        );

    \I__9330\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37147\
        );

    \I__9329\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37140\
        );

    \I__9328\ : InMux
    port map (
            O => \N__37295\,
            I => \N__37140\
        );

    \I__9327\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37140\
        );

    \I__9326\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37137\
        );

    \I__9325\ : Span4Mux_v
    port map (
            O => \N__37290\,
            I => \N__37129\
        );

    \I__9324\ : Span4Mux_h
    port map (
            O => \N__37287\,
            I => \N__37129\
        );

    \I__9323\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37126\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__37281\,
            I => \N__37123\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__37278\,
            I => \N__37118\
        );

    \I__9320\ : Span4Mux_h
    port map (
            O => \N__37273\,
            I => \N__37118\
        );

    \I__9319\ : IoSpan4Mux
    port map (
            O => \N__37270\,
            I => \N__37113\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__37265\,
            I => \N__37113\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__37260\,
            I => \N__37108\
        );

    \I__9316\ : Span4Mux_s3_v
    port map (
            O => \N__37255\,
            I => \N__37108\
        );

    \I__9315\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37105\
        );

    \I__9314\ : InMux
    port map (
            O => \N__37253\,
            I => \N__37098\
        );

    \I__9313\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37098\
        );

    \I__9312\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37098\
        );

    \I__9311\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37093\
        );

    \I__9310\ : InMux
    port map (
            O => \N__37249\,
            I => \N__37093\
        );

    \I__9309\ : InMux
    port map (
            O => \N__37246\,
            I => \N__37090\
        );

    \I__9308\ : CascadeMux
    port map (
            O => \N__37245\,
            I => \N__37085\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__37236\,
            I => \N__37072\
        );

    \I__9306\ : Span4Mux_h
    port map (
            O => \N__37231\,
            I => \N__37061\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__37228\,
            I => \N__37054\
        );

    \I__9304\ : Span4Mux_v
    port map (
            O => \N__37221\,
            I => \N__37054\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__37218\,
            I => \N__37054\
        );

    \I__9302\ : InMux
    port map (
            O => \N__37217\,
            I => \N__37049\
        );

    \I__9301\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37049\
        );

    \I__9300\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37044\
        );

    \I__9299\ : InMux
    port map (
            O => \N__37214\,
            I => \N__37044\
        );

    \I__9298\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37037\
        );

    \I__9297\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37037\
        );

    \I__9296\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37037\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__37206\,
            I => \N__37034\
        );

    \I__9294\ : Span4Mux_h
    port map (
            O => \N__37203\,
            I => \N__37029\
        );

    \I__9293\ : Span4Mux_v
    port map (
            O => \N__37194\,
            I => \N__37029\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__37183\,
            I => \N__37012\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__37180\,
            I => \N__37012\
        );

    \I__9290\ : Span4Mux_h
    port map (
            O => \N__37177\,
            I => \N__37012\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37012\
        );

    \I__9288\ : Span4Mux_v
    port map (
            O => \N__37163\,
            I => \N__37012\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__37154\,
            I => \N__37012\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__37147\,
            I => \N__37012\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__37140\,
            I => \N__37012\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__37137\,
            I => \N__37009\
        );

    \I__9283\ : InMux
    port map (
            O => \N__37136\,
            I => \N__37002\
        );

    \I__9282\ : InMux
    port map (
            O => \N__37135\,
            I => \N__37002\
        );

    \I__9281\ : InMux
    port map (
            O => \N__37134\,
            I => \N__37002\
        );

    \I__9280\ : Span4Mux_h
    port map (
            O => \N__37129\,
            I => \N__36991\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__37126\,
            I => \N__36991\
        );

    \I__9278\ : Span4Mux_h
    port map (
            O => \N__37123\,
            I => \N__36991\
        );

    \I__9277\ : Span4Mux_v
    port map (
            O => \N__37118\,
            I => \N__36991\
        );

    \I__9276\ : Span4Mux_s2_h
    port map (
            O => \N__37113\,
            I => \N__36991\
        );

    \I__9275\ : Span4Mux_h
    port map (
            O => \N__37108\,
            I => \N__36986\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__37105\,
            I => \N__36986\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__37098\,
            I => \N__36983\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__37093\,
            I => \N__36980\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__37090\,
            I => \N__36977\
        );

    \I__9270\ : InMux
    port map (
            O => \N__37089\,
            I => \N__36970\
        );

    \I__9269\ : InMux
    port map (
            O => \N__37088\,
            I => \N__36970\
        );

    \I__9268\ : InMux
    port map (
            O => \N__37085\,
            I => \N__36970\
        );

    \I__9267\ : InMux
    port map (
            O => \N__37084\,
            I => \N__36963\
        );

    \I__9266\ : InMux
    port map (
            O => \N__37083\,
            I => \N__36963\
        );

    \I__9265\ : InMux
    port map (
            O => \N__37082\,
            I => \N__36963\
        );

    \I__9264\ : InMux
    port map (
            O => \N__37081\,
            I => \N__36954\
        );

    \I__9263\ : InMux
    port map (
            O => \N__37080\,
            I => \N__36954\
        );

    \I__9262\ : InMux
    port map (
            O => \N__37079\,
            I => \N__36954\
        );

    \I__9261\ : InMux
    port map (
            O => \N__37078\,
            I => \N__36954\
        );

    \I__9260\ : InMux
    port map (
            O => \N__37077\,
            I => \N__36947\
        );

    \I__9259\ : InMux
    port map (
            O => \N__37076\,
            I => \N__36947\
        );

    \I__9258\ : InMux
    port map (
            O => \N__37075\,
            I => \N__36947\
        );

    \I__9257\ : Span12Mux_s9_h
    port map (
            O => \N__37072\,
            I => \N__36944\
        );

    \I__9256\ : InMux
    port map (
            O => \N__37071\,
            I => \N__36937\
        );

    \I__9255\ : InMux
    port map (
            O => \N__37070\,
            I => \N__36937\
        );

    \I__9254\ : InMux
    port map (
            O => \N__37069\,
            I => \N__36937\
        );

    \I__9253\ : InMux
    port map (
            O => \N__37068\,
            I => \N__36926\
        );

    \I__9252\ : InMux
    port map (
            O => \N__37067\,
            I => \N__36926\
        );

    \I__9251\ : InMux
    port map (
            O => \N__37066\,
            I => \N__36926\
        );

    \I__9250\ : InMux
    port map (
            O => \N__37065\,
            I => \N__36926\
        );

    \I__9249\ : InMux
    port map (
            O => \N__37064\,
            I => \N__36926\
        );

    \I__9248\ : Span4Mux_h
    port map (
            O => \N__37061\,
            I => \N__36919\
        );

    \I__9247\ : Span4Mux_v
    port map (
            O => \N__37054\,
            I => \N__36919\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__37049\,
            I => \N__36919\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__37044\,
            I => \N__36908\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__37037\,
            I => \N__36908\
        );

    \I__9243\ : Span4Mux_v
    port map (
            O => \N__37034\,
            I => \N__36908\
        );

    \I__9242\ : Span4Mux_v
    port map (
            O => \N__37029\,
            I => \N__36908\
        );

    \I__9241\ : Span4Mux_v
    port map (
            O => \N__37012\,
            I => \N__36908\
        );

    \I__9240\ : Span4Mux_h
    port map (
            O => \N__37009\,
            I => \N__36901\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__37002\,
            I => \N__36901\
        );

    \I__9238\ : Span4Mux_v
    port map (
            O => \N__36991\,
            I => \N__36901\
        );

    \I__9237\ : Span4Mux_h
    port map (
            O => \N__36986\,
            I => \N__36890\
        );

    \I__9236\ : Span4Mux_s2_h
    port map (
            O => \N__36983\,
            I => \N__36890\
        );

    \I__9235\ : Span4Mux_v
    port map (
            O => \N__36980\,
            I => \N__36890\
        );

    \I__9234\ : Span4Mux_h
    port map (
            O => \N__36977\,
            I => \N__36890\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__36970\,
            I => \N__36890\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__36963\,
            I => \N__36885\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__36954\,
            I => \N__36885\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__36947\,
            I => instruction_4
        );

    \I__9229\ : Odrv12
    port map (
            O => \N__36944\,
            I => instruction_4
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__36937\,
            I => instruction_4
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__36926\,
            I => instruction_4
        );

    \I__9226\ : Odrv4
    port map (
            O => \N__36919\,
            I => instruction_4
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__36908\,
            I => instruction_4
        );

    \I__9224\ : Odrv4
    port map (
            O => \N__36901\,
            I => instruction_4
        );

    \I__9223\ : Odrv4
    port map (
            O => \N__36890\,
            I => instruction_4
        );

    \I__9222\ : Odrv12
    port map (
            O => \N__36885\,
            I => instruction_4
        );

    \I__9221\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36863\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__36863\,
            I => \N__36860\
        );

    \I__9219\ : Span4Mux_v
    port map (
            O => \N__36860\,
            I => \N__36857\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__36857\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_3\
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__36854\,
            I => \N__36837\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__36853\,
            I => \N__36826\
        );

    \I__9215\ : CascadeMux
    port map (
            O => \N__36852\,
            I => \N__36823\
        );

    \I__9214\ : CascadeMux
    port map (
            O => \N__36851\,
            I => \N__36820\
        );

    \I__9213\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36815\
        );

    \I__9212\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36804\
        );

    \I__9211\ : CascadeMux
    port map (
            O => \N__36848\,
            I => \N__36800\
        );

    \I__9210\ : InMux
    port map (
            O => \N__36847\,
            I => \N__36775\
        );

    \I__9209\ : InMux
    port map (
            O => \N__36846\,
            I => \N__36775\
        );

    \I__9208\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36775\
        );

    \I__9207\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36775\
        );

    \I__9206\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36775\
        );

    \I__9205\ : InMux
    port map (
            O => \N__36842\,
            I => \N__36775\
        );

    \I__9204\ : InMux
    port map (
            O => \N__36841\,
            I => \N__36775\
        );

    \I__9203\ : InMux
    port map (
            O => \N__36840\,
            I => \N__36775\
        );

    \I__9202\ : InMux
    port map (
            O => \N__36837\,
            I => \N__36772\
        );

    \I__9201\ : InMux
    port map (
            O => \N__36836\,
            I => \N__36761\
        );

    \I__9200\ : InMux
    port map (
            O => \N__36835\,
            I => \N__36761\
        );

    \I__9199\ : InMux
    port map (
            O => \N__36834\,
            I => \N__36761\
        );

    \I__9198\ : InMux
    port map (
            O => \N__36833\,
            I => \N__36761\
        );

    \I__9197\ : InMux
    port map (
            O => \N__36832\,
            I => \N__36761\
        );

    \I__9196\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36744\
        );

    \I__9195\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36744\
        );

    \I__9194\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36744\
        );

    \I__9193\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36744\
        );

    \I__9192\ : InMux
    port map (
            O => \N__36823\,
            I => \N__36744\
        );

    \I__9191\ : InMux
    port map (
            O => \N__36820\,
            I => \N__36744\
        );

    \I__9190\ : InMux
    port map (
            O => \N__36819\,
            I => \N__36744\
        );

    \I__9189\ : InMux
    port map (
            O => \N__36818\,
            I => \N__36744\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__36815\,
            I => \N__36733\
        );

    \I__9187\ : InMux
    port map (
            O => \N__36814\,
            I => \N__36716\
        );

    \I__9186\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36716\
        );

    \I__9185\ : InMux
    port map (
            O => \N__36812\,
            I => \N__36716\
        );

    \I__9184\ : InMux
    port map (
            O => \N__36811\,
            I => \N__36716\
        );

    \I__9183\ : InMux
    port map (
            O => \N__36810\,
            I => \N__36716\
        );

    \I__9182\ : InMux
    port map (
            O => \N__36809\,
            I => \N__36716\
        );

    \I__9181\ : InMux
    port map (
            O => \N__36808\,
            I => \N__36716\
        );

    \I__9180\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36716\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__36804\,
            I => \N__36713\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__36803\,
            I => \N__36702\
        );

    \I__9177\ : InMux
    port map (
            O => \N__36800\,
            I => \N__36689\
        );

    \I__9176\ : InMux
    port map (
            O => \N__36799\,
            I => \N__36675\
        );

    \I__9175\ : InMux
    port map (
            O => \N__36798\,
            I => \N__36675\
        );

    \I__9174\ : InMux
    port map (
            O => \N__36797\,
            I => \N__36675\
        );

    \I__9173\ : InMux
    port map (
            O => \N__36796\,
            I => \N__36675\
        );

    \I__9172\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36675\
        );

    \I__9171\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36675\
        );

    \I__9170\ : CascadeMux
    port map (
            O => \N__36793\,
            I => \N__36672\
        );

    \I__9169\ : CascadeMux
    port map (
            O => \N__36792\,
            I => \N__36669\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__36775\,
            I => \N__36652\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__36772\,
            I => \N__36645\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__36761\,
            I => \N__36645\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__36744\,
            I => \N__36645\
        );

    \I__9164\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36628\
        );

    \I__9163\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36628\
        );

    \I__9162\ : InMux
    port map (
            O => \N__36741\,
            I => \N__36628\
        );

    \I__9161\ : InMux
    port map (
            O => \N__36740\,
            I => \N__36628\
        );

    \I__9160\ : InMux
    port map (
            O => \N__36739\,
            I => \N__36628\
        );

    \I__9159\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36628\
        );

    \I__9158\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36628\
        );

    \I__9157\ : InMux
    port map (
            O => \N__36736\,
            I => \N__36628\
        );

    \I__9156\ : Span4Mux_v
    port map (
            O => \N__36733\,
            I => \N__36588\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__36716\,
            I => \N__36588\
        );

    \I__9154\ : Span4Mux_v
    port map (
            O => \N__36713\,
            I => \N__36585\
        );

    \I__9153\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36568\
        );

    \I__9152\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36568\
        );

    \I__9151\ : InMux
    port map (
            O => \N__36710\,
            I => \N__36568\
        );

    \I__9150\ : InMux
    port map (
            O => \N__36709\,
            I => \N__36568\
        );

    \I__9149\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36568\
        );

    \I__9148\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36568\
        );

    \I__9147\ : InMux
    port map (
            O => \N__36706\,
            I => \N__36568\
        );

    \I__9146\ : InMux
    port map (
            O => \N__36705\,
            I => \N__36568\
        );

    \I__9145\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36565\
        );

    \I__9144\ : CascadeMux
    port map (
            O => \N__36701\,
            I => \N__36562\
        );

    \I__9143\ : CascadeMux
    port map (
            O => \N__36700\,
            I => \N__36559\
        );

    \I__9142\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36527\
        );

    \I__9141\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36527\
        );

    \I__9140\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36527\
        );

    \I__9139\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36527\
        );

    \I__9138\ : InMux
    port map (
            O => \N__36695\,
            I => \N__36527\
        );

    \I__9137\ : InMux
    port map (
            O => \N__36694\,
            I => \N__36527\
        );

    \I__9136\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36527\
        );

    \I__9135\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36527\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36519\
        );

    \I__9133\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36516\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__36675\,
            I => \N__36513\
        );

    \I__9131\ : InMux
    port map (
            O => \N__36672\,
            I => \N__36510\
        );

    \I__9130\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36507\
        );

    \I__9129\ : InMux
    port map (
            O => \N__36668\,
            I => \N__36504\
        );

    \I__9128\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36488\
        );

    \I__9127\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36488\
        );

    \I__9126\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36488\
        );

    \I__9125\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36488\
        );

    \I__9124\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36488\
        );

    \I__9123\ : InMux
    port map (
            O => \N__36662\,
            I => \N__36488\
        );

    \I__9122\ : InMux
    port map (
            O => \N__36661\,
            I => \N__36485\
        );

    \I__9121\ : InMux
    port map (
            O => \N__36660\,
            I => \N__36477\
        );

    \I__9120\ : InMux
    port map (
            O => \N__36659\,
            I => \N__36477\
        );

    \I__9119\ : InMux
    port map (
            O => \N__36658\,
            I => \N__36477\
        );

    \I__9118\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36470\
        );

    \I__9117\ : InMux
    port map (
            O => \N__36656\,
            I => \N__36470\
        );

    \I__9116\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36470\
        );

    \I__9115\ : Span4Mux_v
    port map (
            O => \N__36652\,
            I => \N__36467\
        );

    \I__9114\ : Span4Mux_v
    port map (
            O => \N__36645\,
            I => \N__36462\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__36628\,
            I => \N__36462\
        );

    \I__9112\ : CascadeMux
    port map (
            O => \N__36627\,
            I => \N__36459\
        );

    \I__9111\ : CascadeMux
    port map (
            O => \N__36626\,
            I => \N__36456\
        );

    \I__9110\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36450\
        );

    \I__9109\ : InMux
    port map (
            O => \N__36624\,
            I => \N__36450\
        );

    \I__9108\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36447\
        );

    \I__9107\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36430\
        );

    \I__9106\ : InMux
    port map (
            O => \N__36621\,
            I => \N__36430\
        );

    \I__9105\ : InMux
    port map (
            O => \N__36620\,
            I => \N__36430\
        );

    \I__9104\ : InMux
    port map (
            O => \N__36619\,
            I => \N__36430\
        );

    \I__9103\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36430\
        );

    \I__9102\ : InMux
    port map (
            O => \N__36617\,
            I => \N__36430\
        );

    \I__9101\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36430\
        );

    \I__9100\ : InMux
    port map (
            O => \N__36615\,
            I => \N__36430\
        );

    \I__9099\ : InMux
    port map (
            O => \N__36614\,
            I => \N__36415\
        );

    \I__9098\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36415\
        );

    \I__9097\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36415\
        );

    \I__9096\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36415\
        );

    \I__9095\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36415\
        );

    \I__9094\ : InMux
    port map (
            O => \N__36609\,
            I => \N__36415\
        );

    \I__9093\ : InMux
    port map (
            O => \N__36608\,
            I => \N__36415\
        );

    \I__9092\ : CascadeMux
    port map (
            O => \N__36607\,
            I => \N__36407\
        );

    \I__9091\ : CascadeMux
    port map (
            O => \N__36606\,
            I => \N__36400\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__36605\,
            I => \N__36397\
        );

    \I__9089\ : InMux
    port map (
            O => \N__36604\,
            I => \N__36386\
        );

    \I__9088\ : InMux
    port map (
            O => \N__36603\,
            I => \N__36386\
        );

    \I__9087\ : InMux
    port map (
            O => \N__36602\,
            I => \N__36386\
        );

    \I__9086\ : InMux
    port map (
            O => \N__36601\,
            I => \N__36386\
        );

    \I__9085\ : InMux
    port map (
            O => \N__36600\,
            I => \N__36386\
        );

    \I__9084\ : CascadeMux
    port map (
            O => \N__36599\,
            I => \N__36374\
        );

    \I__9083\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36353\
        );

    \I__9082\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36353\
        );

    \I__9081\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36353\
        );

    \I__9080\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36353\
        );

    \I__9079\ : InMux
    port map (
            O => \N__36594\,
            I => \N__36353\
        );

    \I__9078\ : InMux
    port map (
            O => \N__36593\,
            I => \N__36353\
        );

    \I__9077\ : Span4Mux_h
    port map (
            O => \N__36588\,
            I => \N__36344\
        );

    \I__9076\ : Span4Mux_h
    port map (
            O => \N__36585\,
            I => \N__36344\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__36568\,
            I => \N__36344\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__36565\,
            I => \N__36344\
        );

    \I__9073\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36341\
        );

    \I__9072\ : InMux
    port map (
            O => \N__36559\,
            I => \N__36338\
        );

    \I__9071\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36333\
        );

    \I__9070\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36333\
        );

    \I__9069\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36316\
        );

    \I__9068\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36316\
        );

    \I__9067\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36316\
        );

    \I__9066\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36316\
        );

    \I__9065\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36316\
        );

    \I__9064\ : InMux
    port map (
            O => \N__36551\,
            I => \N__36316\
        );

    \I__9063\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36316\
        );

    \I__9062\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36316\
        );

    \I__9061\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36298\
        );

    \I__9060\ : InMux
    port map (
            O => \N__36547\,
            I => \N__36298\
        );

    \I__9059\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36298\
        );

    \I__9058\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36298\
        );

    \I__9057\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36298\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__36527\,
            I => \N__36295\
        );

    \I__9055\ : InMux
    port map (
            O => \N__36526\,
            I => \N__36288\
        );

    \I__9054\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36288\
        );

    \I__9053\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36288\
        );

    \I__9052\ : CascadeMux
    port map (
            O => \N__36523\,
            I => \N__36285\
        );

    \I__9051\ : CascadeMux
    port map (
            O => \N__36522\,
            I => \N__36276\
        );

    \I__9050\ : Span4Mux_v
    port map (
            O => \N__36519\,
            I => \N__36263\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__36516\,
            I => \N__36263\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__36513\,
            I => \N__36263\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__36510\,
            I => \N__36263\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__36507\,
            I => \N__36263\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__36504\,
            I => \N__36263\
        );

    \I__9044\ : InMux
    port map (
            O => \N__36503\,
            I => \N__36258\
        );

    \I__9043\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36258\
        );

    \I__9042\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36255\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__36488\,
            I => \N__36252\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__36485\,
            I => \N__36249\
        );

    \I__9039\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36246\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__36477\,
            I => \N__36237\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__36470\,
            I => \N__36237\
        );

    \I__9036\ : Span4Mux_s0_h
    port map (
            O => \N__36467\,
            I => \N__36237\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__36462\,
            I => \N__36237\
        );

    \I__9034\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36234\
        );

    \I__9033\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36231\
        );

    \I__9032\ : InMux
    port map (
            O => \N__36455\,
            I => \N__36228\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__36450\,
            I => \N__36223\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__36447\,
            I => \N__36223\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__36430\,
            I => \N__36218\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__36415\,
            I => \N__36218\
        );

    \I__9027\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36207\
        );

    \I__9026\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36207\
        );

    \I__9025\ : InMux
    port map (
            O => \N__36412\,
            I => \N__36207\
        );

    \I__9024\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36207\
        );

    \I__9023\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36207\
        );

    \I__9022\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36204\
        );

    \I__9021\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36168\
        );

    \I__9020\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36168\
        );

    \I__9019\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36168\
        );

    \I__9018\ : InMux
    port map (
            O => \N__36403\,
            I => \N__36168\
        );

    \I__9017\ : InMux
    port map (
            O => \N__36400\,
            I => \N__36168\
        );

    \I__9016\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36168\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__36386\,
            I => \N__36165\
        );

    \I__9014\ : InMux
    port map (
            O => \N__36385\,
            I => \N__36148\
        );

    \I__9013\ : InMux
    port map (
            O => \N__36384\,
            I => \N__36148\
        );

    \I__9012\ : InMux
    port map (
            O => \N__36383\,
            I => \N__36148\
        );

    \I__9011\ : InMux
    port map (
            O => \N__36382\,
            I => \N__36148\
        );

    \I__9010\ : InMux
    port map (
            O => \N__36381\,
            I => \N__36148\
        );

    \I__9009\ : InMux
    port map (
            O => \N__36380\,
            I => \N__36148\
        );

    \I__9008\ : InMux
    port map (
            O => \N__36379\,
            I => \N__36148\
        );

    \I__9007\ : InMux
    port map (
            O => \N__36378\,
            I => \N__36148\
        );

    \I__9006\ : InMux
    port map (
            O => \N__36377\,
            I => \N__36145\
        );

    \I__9005\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36134\
        );

    \I__9004\ : InMux
    port map (
            O => \N__36373\,
            I => \N__36117\
        );

    \I__9003\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36117\
        );

    \I__9002\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36117\
        );

    \I__9001\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36117\
        );

    \I__9000\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36117\
        );

    \I__8999\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36117\
        );

    \I__8998\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36117\
        );

    \I__8997\ : InMux
    port map (
            O => \N__36366\,
            I => \N__36117\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__36353\,
            I => \N__36112\
        );

    \I__8995\ : Span4Mux_v
    port map (
            O => \N__36344\,
            I => \N__36112\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__36341\,
            I => \N__36103\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__36338\,
            I => \N__36103\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__36333\,
            I => \N__36103\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__36316\,
            I => \N__36103\
        );

    \I__8990\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36095\
        );

    \I__8989\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36082\
        );

    \I__8988\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36082\
        );

    \I__8987\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36082\
        );

    \I__8986\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36082\
        );

    \I__8985\ : InMux
    port map (
            O => \N__36310\,
            I => \N__36082\
        );

    \I__8984\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36082\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__36298\,
            I => \N__36079\
        );

    \I__8982\ : Span4Mux_v
    port map (
            O => \N__36295\,
            I => \N__36074\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__36288\,
            I => \N__36074\
        );

    \I__8980\ : InMux
    port map (
            O => \N__36285\,
            I => \N__36071\
        );

    \I__8979\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36058\
        );

    \I__8978\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36058\
        );

    \I__8977\ : InMux
    port map (
            O => \N__36282\,
            I => \N__36058\
        );

    \I__8976\ : InMux
    port map (
            O => \N__36281\,
            I => \N__36058\
        );

    \I__8975\ : InMux
    port map (
            O => \N__36280\,
            I => \N__36058\
        );

    \I__8974\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36058\
        );

    \I__8973\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36055\
        );

    \I__8972\ : Span4Mux_h
    port map (
            O => \N__36263\,
            I => \N__36052\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__36258\,
            I => \N__36035\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__36255\,
            I => \N__36035\
        );

    \I__8969\ : Span4Mux_v
    port map (
            O => \N__36252\,
            I => \N__36035\
        );

    \I__8968\ : Span4Mux_s3_h
    port map (
            O => \N__36249\,
            I => \N__36035\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__36246\,
            I => \N__36035\
        );

    \I__8966\ : Span4Mux_h
    port map (
            O => \N__36237\,
            I => \N__36035\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__36234\,
            I => \N__36035\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__36231\,
            I => \N__36029\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__36228\,
            I => \N__36029\
        );

    \I__8962\ : Span4Mux_s3_v
    port map (
            O => \N__36223\,
            I => \N__36024\
        );

    \I__8961\ : Span4Mux_h
    port map (
            O => \N__36218\,
            I => \N__36024\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__36207\,
            I => \N__36019\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__36204\,
            I => \N__36019\
        );

    \I__8958\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36002\
        );

    \I__8957\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36002\
        );

    \I__8956\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36002\
        );

    \I__8955\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36002\
        );

    \I__8954\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36002\
        );

    \I__8953\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36002\
        );

    \I__8952\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36002\
        );

    \I__8951\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36002\
        );

    \I__8950\ : CascadeMux
    port map (
            O => \N__36195\,
            I => \N__35999\
        );

    \I__8949\ : CascadeMux
    port map (
            O => \N__36194\,
            I => \N__35996\
        );

    \I__8948\ : InMux
    port map (
            O => \N__36193\,
            I => \N__35952\
        );

    \I__8947\ : InMux
    port map (
            O => \N__36192\,
            I => \N__35952\
        );

    \I__8946\ : InMux
    port map (
            O => \N__36191\,
            I => \N__35952\
        );

    \I__8945\ : InMux
    port map (
            O => \N__36190\,
            I => \N__35952\
        );

    \I__8944\ : InMux
    port map (
            O => \N__36189\,
            I => \N__35952\
        );

    \I__8943\ : InMux
    port map (
            O => \N__36188\,
            I => \N__35952\
        );

    \I__8942\ : InMux
    port map (
            O => \N__36187\,
            I => \N__35952\
        );

    \I__8941\ : InMux
    port map (
            O => \N__36186\,
            I => \N__35952\
        );

    \I__8940\ : InMux
    port map (
            O => \N__36185\,
            I => \N__35941\
        );

    \I__8939\ : InMux
    port map (
            O => \N__36184\,
            I => \N__35941\
        );

    \I__8938\ : InMux
    port map (
            O => \N__36183\,
            I => \N__35941\
        );

    \I__8937\ : InMux
    port map (
            O => \N__36182\,
            I => \N__35941\
        );

    \I__8936\ : InMux
    port map (
            O => \N__36181\,
            I => \N__35941\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__36168\,
            I => \N__35934\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__36165\,
            I => \N__35934\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__36148\,
            I => \N__35934\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__36145\,
            I => \N__35931\
        );

    \I__8931\ : InMux
    port map (
            O => \N__36144\,
            I => \N__35926\
        );

    \I__8930\ : InMux
    port map (
            O => \N__36143\,
            I => \N__35926\
        );

    \I__8929\ : InMux
    port map (
            O => \N__36142\,
            I => \N__35913\
        );

    \I__8928\ : InMux
    port map (
            O => \N__36141\,
            I => \N__35913\
        );

    \I__8927\ : InMux
    port map (
            O => \N__36140\,
            I => \N__35913\
        );

    \I__8926\ : InMux
    port map (
            O => \N__36139\,
            I => \N__35913\
        );

    \I__8925\ : InMux
    port map (
            O => \N__36138\,
            I => \N__35913\
        );

    \I__8924\ : InMux
    port map (
            O => \N__36137\,
            I => \N__35913\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__36134\,
            I => \N__35910\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__36117\,
            I => \N__35907\
        );

    \I__8921\ : Span4Mux_h
    port map (
            O => \N__36112\,
            I => \N__35902\
        );

    \I__8920\ : Span4Mux_v
    port map (
            O => \N__36103\,
            I => \N__35902\
        );

    \I__8919\ : InMux
    port map (
            O => \N__36102\,
            I => \N__35899\
        );

    \I__8918\ : InMux
    port map (
            O => \N__36101\,
            I => \N__35896\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__36100\,
            I => \N__35893\
        );

    \I__8916\ : CascadeMux
    port map (
            O => \N__36099\,
            I => \N__35890\
        );

    \I__8915\ : CascadeMux
    port map (
            O => \N__36098\,
            I => \N__35887\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__36095\,
            I => \N__35871\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__36082\,
            I => \N__35871\
        );

    \I__8912\ : Span4Mux_s3_h
    port map (
            O => \N__36079\,
            I => \N__35862\
        );

    \I__8911\ : Span4Mux_h
    port map (
            O => \N__36074\,
            I => \N__35862\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__35862\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__36058\,
            I => \N__35862\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__36055\,
            I => \N__35854\
        );

    \I__8907\ : Span4Mux_h
    port map (
            O => \N__36052\,
            I => \N__35854\
        );

    \I__8906\ : InMux
    port map (
            O => \N__36051\,
            I => \N__35849\
        );

    \I__8905\ : InMux
    port map (
            O => \N__36050\,
            I => \N__35849\
        );

    \I__8904\ : Span4Mux_h
    port map (
            O => \N__36035\,
            I => \N__35840\
        );

    \I__8903\ : InMux
    port map (
            O => \N__36034\,
            I => \N__35837\
        );

    \I__8902\ : Span4Mux_s3_v
    port map (
            O => \N__36029\,
            I => \N__35832\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__36024\,
            I => \N__35832\
        );

    \I__8900\ : Span4Mux_h
    port map (
            O => \N__36019\,
            I => \N__35827\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__36002\,
            I => \N__35827\
        );

    \I__8898\ : InMux
    port map (
            O => \N__35999\,
            I => \N__35822\
        );

    \I__8897\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35822\
        );

    \I__8896\ : InMux
    port map (
            O => \N__35995\,
            I => \N__35809\
        );

    \I__8895\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35809\
        );

    \I__8894\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35809\
        );

    \I__8893\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35809\
        );

    \I__8892\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35809\
        );

    \I__8891\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35809\
        );

    \I__8890\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35798\
        );

    \I__8889\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35798\
        );

    \I__8888\ : InMux
    port map (
            O => \N__35987\,
            I => \N__35798\
        );

    \I__8887\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35798\
        );

    \I__8886\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35798\
        );

    \I__8885\ : InMux
    port map (
            O => \N__35984\,
            I => \N__35791\
        );

    \I__8884\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35791\
        );

    \I__8883\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35791\
        );

    \I__8882\ : InMux
    port map (
            O => \N__35981\,
            I => \N__35778\
        );

    \I__8881\ : InMux
    port map (
            O => \N__35980\,
            I => \N__35778\
        );

    \I__8880\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35778\
        );

    \I__8879\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35778\
        );

    \I__8878\ : InMux
    port map (
            O => \N__35977\,
            I => \N__35778\
        );

    \I__8877\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35778\
        );

    \I__8876\ : InMux
    port map (
            O => \N__35975\,
            I => \N__35763\
        );

    \I__8875\ : InMux
    port map (
            O => \N__35974\,
            I => \N__35763\
        );

    \I__8874\ : InMux
    port map (
            O => \N__35973\,
            I => \N__35763\
        );

    \I__8873\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35763\
        );

    \I__8872\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35763\
        );

    \I__8871\ : InMux
    port map (
            O => \N__35970\,
            I => \N__35763\
        );

    \I__8870\ : InMux
    port map (
            O => \N__35969\,
            I => \N__35763\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__35952\,
            I => \N__35758\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__35941\,
            I => \N__35758\
        );

    \I__8867\ : Span4Mux_h
    port map (
            O => \N__35934\,
            I => \N__35755\
        );

    \I__8866\ : Span4Mux_v
    port map (
            O => \N__35931\,
            I => \N__35750\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__35926\,
            I => \N__35750\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__35913\,
            I => \N__35747\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__35910\,
            I => \N__35742\
        );

    \I__8862\ : Span4Mux_v
    port map (
            O => \N__35907\,
            I => \N__35737\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__35902\,
            I => \N__35737\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__35899\,
            I => \N__35732\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35732\
        );

    \I__8858\ : InMux
    port map (
            O => \N__35893\,
            I => \N__35727\
        );

    \I__8857\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35724\
        );

    \I__8856\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35715\
        );

    \I__8855\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35715\
        );

    \I__8854\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35715\
        );

    \I__8853\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35715\
        );

    \I__8852\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35698\
        );

    \I__8851\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35698\
        );

    \I__8850\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35698\
        );

    \I__8849\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35698\
        );

    \I__8848\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35698\
        );

    \I__8847\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35698\
        );

    \I__8846\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35698\
        );

    \I__8845\ : InMux
    port map (
            O => \N__35876\,
            I => \N__35698\
        );

    \I__8844\ : Span4Mux_s2_v
    port map (
            O => \N__35871\,
            I => \N__35693\
        );

    \I__8843\ : Span4Mux_v
    port map (
            O => \N__35862\,
            I => \N__35693\
        );

    \I__8842\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35686\
        );

    \I__8841\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35686\
        );

    \I__8840\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35686\
        );

    \I__8839\ : Sp12to4
    port map (
            O => \N__35854\,
            I => \N__35681\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__35849\,
            I => \N__35681\
        );

    \I__8837\ : InMux
    port map (
            O => \N__35848\,
            I => \N__35668\
        );

    \I__8836\ : InMux
    port map (
            O => \N__35847\,
            I => \N__35668\
        );

    \I__8835\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35668\
        );

    \I__8834\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35668\
        );

    \I__8833\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35668\
        );

    \I__8832\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35668\
        );

    \I__8831\ : Sp12to4
    port map (
            O => \N__35840\,
            I => \N__35663\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__35837\,
            I => \N__35663\
        );

    \I__8829\ : Span4Mux_v
    port map (
            O => \N__35832\,
            I => \N__35658\
        );

    \I__8828\ : Span4Mux_s3_h
    port map (
            O => \N__35827\,
            I => \N__35658\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__35822\,
            I => \N__35649\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__35809\,
            I => \N__35649\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__35798\,
            I => \N__35649\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__35791\,
            I => \N__35649\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35644\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__35763\,
            I => \N__35644\
        );

    \I__8821\ : Span4Mux_h
    port map (
            O => \N__35758\,
            I => \N__35637\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__35755\,
            I => \N__35637\
        );

    \I__8819\ : Span4Mux_v
    port map (
            O => \N__35750\,
            I => \N__35637\
        );

    \I__8818\ : Span4Mux_h
    port map (
            O => \N__35747\,
            I => \N__35634\
        );

    \I__8817\ : InMux
    port map (
            O => \N__35746\,
            I => \N__35629\
        );

    \I__8816\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35629\
        );

    \I__8815\ : Span4Mux_h
    port map (
            O => \N__35742\,
            I => \N__35622\
        );

    \I__8814\ : Span4Mux_v
    port map (
            O => \N__35737\,
            I => \N__35622\
        );

    \I__8813\ : Span4Mux_s2_v
    port map (
            O => \N__35732\,
            I => \N__35622\
        );

    \I__8812\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35617\
        );

    \I__8811\ : InMux
    port map (
            O => \N__35730\,
            I => \N__35617\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__35727\,
            I => \N__35600\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__35724\,
            I => \N__35600\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__35715\,
            I => \N__35600\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__35698\,
            I => \N__35600\
        );

    \I__8806\ : Sp12to4
    port map (
            O => \N__35693\,
            I => \N__35600\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__35686\,
            I => \N__35600\
        );

    \I__8804\ : Span12Mux_v
    port map (
            O => \N__35681\,
            I => \N__35600\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__35668\,
            I => \N__35600\
        );

    \I__8802\ : Span12Mux_s8_v
    port map (
            O => \N__35663\,
            I => \N__35593\
        );

    \I__8801\ : Sp12to4
    port map (
            O => \N__35658\,
            I => \N__35593\
        );

    \I__8800\ : Span12Mux_s8_h
    port map (
            O => \N__35649\,
            I => \N__35593\
        );

    \I__8799\ : Span4Mux_h
    port map (
            O => \N__35644\,
            I => \N__35588\
        );

    \I__8798\ : Span4Mux_h
    port map (
            O => \N__35637\,
            I => \N__35588\
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__35634\,
            I => \processor_zipi8.alu_mux_sel_1\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__35629\,
            I => \processor_zipi8.alu_mux_sel_1\
        );

    \I__8795\ : Odrv4
    port map (
            O => \N__35622\,
            I => \processor_zipi8.alu_mux_sel_1\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__35617\,
            I => \processor_zipi8.alu_mux_sel_1\
        );

    \I__8793\ : Odrv12
    port map (
            O => \N__35600\,
            I => \processor_zipi8.alu_mux_sel_1\
        );

    \I__8792\ : Odrv12
    port map (
            O => \N__35593\,
            I => \processor_zipi8.alu_mux_sel_1\
        );

    \I__8791\ : Odrv4
    port map (
            O => \N__35588\,
            I => \processor_zipi8.alu_mux_sel_1\
        );

    \I__8790\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35570\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__35570\,
            I => \N__35564\
        );

    \I__8788\ : CascadeMux
    port map (
            O => \N__35569\,
            I => \N__35561\
        );

    \I__8787\ : CascadeMux
    port map (
            O => \N__35568\,
            I => \N__35553\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__35567\,
            I => \N__35550\
        );

    \I__8785\ : Span4Mux_v
    port map (
            O => \N__35564\,
            I => \N__35542\
        );

    \I__8784\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35539\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__35560\,
            I => \N__35536\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__35559\,
            I => \N__35532\
        );

    \I__8781\ : CascadeMux
    port map (
            O => \N__35558\,
            I => \N__35527\
        );

    \I__8780\ : CascadeMux
    port map (
            O => \N__35557\,
            I => \N__35524\
        );

    \I__8779\ : CascadeMux
    port map (
            O => \N__35556\,
            I => \N__35518\
        );

    \I__8778\ : InMux
    port map (
            O => \N__35553\,
            I => \N__35515\
        );

    \I__8777\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35512\
        );

    \I__8776\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35508\
        );

    \I__8775\ : CascadeMux
    port map (
            O => \N__35548\,
            I => \N__35505\
        );

    \I__8774\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35502\
        );

    \I__8773\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35499\
        );

    \I__8772\ : InMux
    port map (
            O => \N__35545\,
            I => \N__35495\
        );

    \I__8771\ : Span4Mux_s2_h
    port map (
            O => \N__35542\,
            I => \N__35489\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__35539\,
            I => \N__35489\
        );

    \I__8769\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35486\
        );

    \I__8768\ : CascadeMux
    port map (
            O => \N__35535\,
            I => \N__35482\
        );

    \I__8767\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35479\
        );

    \I__8766\ : InMux
    port map (
            O => \N__35531\,
            I => \N__35476\
        );

    \I__8765\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35473\
        );

    \I__8764\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35469\
        );

    \I__8763\ : InMux
    port map (
            O => \N__35524\,
            I => \N__35466\
        );

    \I__8762\ : InMux
    port map (
            O => \N__35523\,
            I => \N__35463\
        );

    \I__8761\ : InMux
    port map (
            O => \N__35522\,
            I => \N__35460\
        );

    \I__8760\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35457\
        );

    \I__8759\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35454\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__35515\,
            I => \N__35449\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N__35449\
        );

    \I__8756\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35446\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35443\
        );

    \I__8754\ : InMux
    port map (
            O => \N__35505\,
            I => \N__35440\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__35502\,
            I => \N__35435\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__35499\,
            I => \N__35435\
        );

    \I__8751\ : InMux
    port map (
            O => \N__35498\,
            I => \N__35432\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__35495\,
            I => \N__35429\
        );

    \I__8749\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35423\
        );

    \I__8748\ : Span4Mux_v
    port map (
            O => \N__35489\,
            I => \N__35418\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__35486\,
            I => \N__35418\
        );

    \I__8746\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35415\
        );

    \I__8745\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35410\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__35479\,
            I => \N__35405\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__35476\,
            I => \N__35405\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__35473\,
            I => \N__35402\
        );

    \I__8741\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35399\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__35469\,
            I => \N__35396\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__35466\,
            I => \N__35393\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__35463\,
            I => \N__35382\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__35460\,
            I => \N__35382\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__35457\,
            I => \N__35382\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__35454\,
            I => \N__35382\
        );

    \I__8734\ : Span4Mux_s2_v
    port map (
            O => \N__35449\,
            I => \N__35382\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__35446\,
            I => \N__35377\
        );

    \I__8732\ : Span4Mux_v
    port map (
            O => \N__35443\,
            I => \N__35377\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__35440\,
            I => \N__35372\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__35435\,
            I => \N__35372\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__35432\,
            I => \N__35367\
        );

    \I__8728\ : Span4Mux_s1_h
    port map (
            O => \N__35429\,
            I => \N__35367\
        );

    \I__8727\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35364\
        );

    \I__8726\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35360\
        );

    \I__8725\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35357\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__35423\,
            I => \N__35354\
        );

    \I__8723\ : Span4Mux_v
    port map (
            O => \N__35418\,
            I => \N__35351\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__35415\,
            I => \N__35348\
        );

    \I__8721\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35344\
        );

    \I__8720\ : CascadeMux
    port map (
            O => \N__35413\,
            I => \N__35341\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__35410\,
            I => \N__35333\
        );

    \I__8718\ : Span4Mux_s1_h
    port map (
            O => \N__35405\,
            I => \N__35333\
        );

    \I__8717\ : Span4Mux_v
    port map (
            O => \N__35402\,
            I => \N__35333\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__35399\,
            I => \N__35328\
        );

    \I__8715\ : Span4Mux_s1_h
    port map (
            O => \N__35396\,
            I => \N__35328\
        );

    \I__8714\ : Span4Mux_s3_h
    port map (
            O => \N__35393\,
            I => \N__35319\
        );

    \I__8713\ : Span4Mux_v
    port map (
            O => \N__35382\,
            I => \N__35319\
        );

    \I__8712\ : Span4Mux_v
    port map (
            O => \N__35377\,
            I => \N__35319\
        );

    \I__8711\ : Span4Mux_v
    port map (
            O => \N__35372\,
            I => \N__35319\
        );

    \I__8710\ : Sp12to4
    port map (
            O => \N__35367\,
            I => \N__35314\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__35364\,
            I => \N__35314\
        );

    \I__8708\ : InMux
    port map (
            O => \N__35363\,
            I => \N__35311\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__35360\,
            I => \N__35306\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__35357\,
            I => \N__35306\
        );

    \I__8705\ : Span4Mux_v
    port map (
            O => \N__35354\,
            I => \N__35303\
        );

    \I__8704\ : Span4Mux_h
    port map (
            O => \N__35351\,
            I => \N__35298\
        );

    \I__8703\ : Span4Mux_s1_h
    port map (
            O => \N__35348\,
            I => \N__35298\
        );

    \I__8702\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35294\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__35344\,
            I => \N__35291\
        );

    \I__8700\ : InMux
    port map (
            O => \N__35341\,
            I => \N__35288\
        );

    \I__8699\ : InMux
    port map (
            O => \N__35340\,
            I => \N__35285\
        );

    \I__8698\ : Span4Mux_h
    port map (
            O => \N__35333\,
            I => \N__35280\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__35328\,
            I => \N__35280\
        );

    \I__8696\ : Sp12to4
    port map (
            O => \N__35319\,
            I => \N__35275\
        );

    \I__8695\ : Span12Mux_s9_v
    port map (
            O => \N__35314\,
            I => \N__35275\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__35311\,
            I => \N__35268\
        );

    \I__8693\ : Span4Mux_v
    port map (
            O => \N__35306\,
            I => \N__35268\
        );

    \I__8692\ : Span4Mux_h
    port map (
            O => \N__35303\,
            I => \N__35268\
        );

    \I__8691\ : Span4Mux_h
    port map (
            O => \N__35298\,
            I => \N__35265\
        );

    \I__8690\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35262\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__35294\,
            I => \N__35255\
        );

    \I__8688\ : Span12Mux_s6_h
    port map (
            O => \N__35291\,
            I => \N__35255\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__35288\,
            I => \N__35255\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__35285\,
            I => \processor_zipi8.arith_logical_result_4\
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__35280\,
            I => \processor_zipi8.arith_logical_result_4\
        );

    \I__8684\ : Odrv12
    port map (
            O => \N__35275\,
            I => \processor_zipi8.arith_logical_result_4\
        );

    \I__8683\ : Odrv4
    port map (
            O => \N__35268\,
            I => \processor_zipi8.arith_logical_result_4\
        );

    \I__8682\ : Odrv4
    port map (
            O => \N__35265\,
            I => \processor_zipi8.arith_logical_result_4\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__35262\,
            I => \processor_zipi8.arith_logical_result_4\
        );

    \I__8680\ : Odrv12
    port map (
            O => \N__35255\,
            I => \processor_zipi8.arith_logical_result_4\
        );

    \I__8679\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35237\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__35237\,
            I => \N__35225\
        );

    \I__8677\ : CascadeMux
    port map (
            O => \N__35236\,
            I => \N__35222\
        );

    \I__8676\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35215\
        );

    \I__8675\ : CascadeMux
    port map (
            O => \N__35234\,
            I => \N__35212\
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__35233\,
            I => \N__35208\
        );

    \I__8673\ : CascadeMux
    port map (
            O => \N__35232\,
            I => \N__35205\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__35231\,
            I => \N__35200\
        );

    \I__8671\ : CascadeMux
    port map (
            O => \N__35230\,
            I => \N__35197\
        );

    \I__8670\ : CascadeMux
    port map (
            O => \N__35229\,
            I => \N__35194\
        );

    \I__8669\ : InMux
    port map (
            O => \N__35228\,
            I => \N__35186\
        );

    \I__8668\ : Span4Mux_v
    port map (
            O => \N__35225\,
            I => \N__35183\
        );

    \I__8667\ : InMux
    port map (
            O => \N__35222\,
            I => \N__35180\
        );

    \I__8666\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35177\
        );

    \I__8665\ : InMux
    port map (
            O => \N__35220\,
            I => \N__35174\
        );

    \I__8664\ : CascadeMux
    port map (
            O => \N__35219\,
            I => \N__35171\
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__35218\,
            I => \N__35166\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__35215\,
            I => \N__35163\
        );

    \I__8661\ : InMux
    port map (
            O => \N__35212\,
            I => \N__35160\
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__35211\,
            I => \N__35157\
        );

    \I__8659\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35152\
        );

    \I__8658\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35149\
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__35204\,
            I => \N__35146\
        );

    \I__8656\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35142\
        );

    \I__8655\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35139\
        );

    \I__8654\ : InMux
    port map (
            O => \N__35197\,
            I => \N__35136\
        );

    \I__8653\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35133\
        );

    \I__8652\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35130\
        );

    \I__8651\ : CascadeMux
    port map (
            O => \N__35192\,
            I => \N__35127\
        );

    \I__8650\ : CascadeMux
    port map (
            O => \N__35191\,
            I => \N__35124\
        );

    \I__8649\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35120\
        );

    \I__8648\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35117\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__35186\,
            I => \N__35114\
        );

    \I__8646\ : IoSpan4Mux
    port map (
            O => \N__35183\,
            I => \N__35107\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__35107\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35107\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__35174\,
            I => \N__35104\
        );

    \I__8642\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35101\
        );

    \I__8641\ : InMux
    port map (
            O => \N__35170\,
            I => \N__35098\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__35169\,
            I => \N__35094\
        );

    \I__8639\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35090\
        );

    \I__8638\ : Span4Mux_v
    port map (
            O => \N__35163\,
            I => \N__35085\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__35160\,
            I => \N__35085\
        );

    \I__8636\ : InMux
    port map (
            O => \N__35157\,
            I => \N__35082\
        );

    \I__8635\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35079\
        );

    \I__8634\ : InMux
    port map (
            O => \N__35155\,
            I => \N__35076\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__35152\,
            I => \N__35073\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__35149\,
            I => \N__35070\
        );

    \I__8631\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35067\
        );

    \I__8630\ : InMux
    port map (
            O => \N__35145\,
            I => \N__35064\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__35142\,
            I => \N__35057\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__35139\,
            I => \N__35057\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__35136\,
            I => \N__35057\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__35133\,
            I => \N__35054\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__35130\,
            I => \N__35051\
        );

    \I__8624\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35048\
        );

    \I__8623\ : InMux
    port map (
            O => \N__35124\,
            I => \N__35045\
        );

    \I__8622\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35042\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__35120\,
            I => \N__35039\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__35117\,
            I => \N__35032\
        );

    \I__8619\ : Span4Mux_v
    port map (
            O => \N__35114\,
            I => \N__35032\
        );

    \I__8618\ : Span4Mux_s2_h
    port map (
            O => \N__35107\,
            I => \N__35032\
        );

    \I__8617\ : Span4Mux_v
    port map (
            O => \N__35104\,
            I => \N__35029\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__35101\,
            I => \N__35024\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__35098\,
            I => \N__35024\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__35097\,
            I => \N__35021\
        );

    \I__8613\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35018\
        );

    \I__8612\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35015\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__35090\,
            I => \N__35008\
        );

    \I__8610\ : Span4Mux_h
    port map (
            O => \N__35085\,
            I => \N__35008\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__35082\,
            I => \N__35008\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__35079\,
            I => \N__35001\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35001\
        );

    \I__8606\ : Span4Mux_s1_h
    port map (
            O => \N__35073\,
            I => \N__34996\
        );

    \I__8605\ : Span4Mux_v
    port map (
            O => \N__35070\,
            I => \N__34996\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__35067\,
            I => \N__34989\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__35064\,
            I => \N__34989\
        );

    \I__8602\ : Span4Mux_s3_v
    port map (
            O => \N__35057\,
            I => \N__34989\
        );

    \I__8601\ : Span4Mux_v
    port map (
            O => \N__35054\,
            I => \N__34986\
        );

    \I__8600\ : Span4Mux_s2_v
    port map (
            O => \N__35051\,
            I => \N__34979\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__35048\,
            I => \N__34979\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__35045\,
            I => \N__34979\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__35042\,
            I => \N__34968\
        );

    \I__8596\ : Span4Mux_v
    port map (
            O => \N__35039\,
            I => \N__34968\
        );

    \I__8595\ : Span4Mux_v
    port map (
            O => \N__35032\,
            I => \N__34968\
        );

    \I__8594\ : Span4Mux_s2_h
    port map (
            O => \N__35029\,
            I => \N__34968\
        );

    \I__8593\ : Span4Mux_s2_h
    port map (
            O => \N__35024\,
            I => \N__34968\
        );

    \I__8592\ : InMux
    port map (
            O => \N__35021\,
            I => \N__34965\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__35018\,
            I => \N__34960\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__35015\,
            I => \N__34960\
        );

    \I__8589\ : Span4Mux_h
    port map (
            O => \N__35008\,
            I => \N__34957\
        );

    \I__8588\ : InMux
    port map (
            O => \N__35007\,
            I => \N__34954\
        );

    \I__8587\ : InMux
    port map (
            O => \N__35006\,
            I => \N__34951\
        );

    \I__8586\ : Span12Mux_s8_v
    port map (
            O => \N__35001\,
            I => \N__34948\
        );

    \I__8585\ : Span4Mux_h
    port map (
            O => \N__34996\,
            I => \N__34945\
        );

    \I__8584\ : Span4Mux_v
    port map (
            O => \N__34989\,
            I => \N__34940\
        );

    \I__8583\ : Span4Mux_v
    port map (
            O => \N__34986\,
            I => \N__34940\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__34979\,
            I => \N__34935\
        );

    \I__8581\ : Span4Mux_h
    port map (
            O => \N__34968\,
            I => \N__34935\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__34965\,
            I => \N__34926\
        );

    \I__8579\ : Span12Mux_s6_h
    port map (
            O => \N__34960\,
            I => \N__34926\
        );

    \I__8578\ : Sp12to4
    port map (
            O => \N__34957\,
            I => \N__34926\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__34954\,
            I => \N__34926\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__34951\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\
        );

    \I__8575\ : Odrv12
    port map (
            O => \N__34948\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__34945\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__34940\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\
        );

    \I__8572\ : Odrv4
    port map (
            O => \N__34935\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\
        );

    \I__8571\ : Odrv12
    port map (
            O => \N__34926\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\
        );

    \I__8570\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34892\
        );

    \I__8569\ : InMux
    port map (
            O => \N__34912\,
            I => \N__34892\
        );

    \I__8568\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34892\
        );

    \I__8567\ : InMux
    port map (
            O => \N__34910\,
            I => \N__34892\
        );

    \I__8566\ : InMux
    port map (
            O => \N__34909\,
            I => \N__34892\
        );

    \I__8565\ : InMux
    port map (
            O => \N__34908\,
            I => \N__34892\
        );

    \I__8564\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34892\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__34892\,
            I => \N__34877\
        );

    \I__8562\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34862\
        );

    \I__8561\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34862\
        );

    \I__8560\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34862\
        );

    \I__8559\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34862\
        );

    \I__8558\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34862\
        );

    \I__8557\ : InMux
    port map (
            O => \N__34886\,
            I => \N__34862\
        );

    \I__8556\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34862\
        );

    \I__8555\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34859\
        );

    \I__8554\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34852\
        );

    \I__8553\ : InMux
    port map (
            O => \N__34882\,
            I => \N__34852\
        );

    \I__8552\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34852\
        );

    \I__8551\ : CascadeMux
    port map (
            O => \N__34880\,
            I => \N__34847\
        );

    \I__8550\ : Span4Mux_v
    port map (
            O => \N__34877\,
            I => \N__34786\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__34862\,
            I => \N__34786\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__34859\,
            I => \N__34786\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__34852\,
            I => \N__34783\
        );

    \I__8546\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34766\
        );

    \I__8545\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34766\
        );

    \I__8544\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34766\
        );

    \I__8543\ : InMux
    port map (
            O => \N__34846\,
            I => \N__34766\
        );

    \I__8542\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34766\
        );

    \I__8541\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34766\
        );

    \I__8540\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34766\
        );

    \I__8539\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34766\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__34841\,
            I => \N__34761\
        );

    \I__8537\ : CascadeMux
    port map (
            O => \N__34840\,
            I => \N__34757\
        );

    \I__8536\ : CascadeMux
    port map (
            O => \N__34839\,
            I => \N__34748\
        );

    \I__8535\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34727\
        );

    \I__8534\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34727\
        );

    \I__8533\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34727\
        );

    \I__8532\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34727\
        );

    \I__8531\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34727\
        );

    \I__8530\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34727\
        );

    \I__8529\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34727\
        );

    \I__8528\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34723\
        );

    \I__8527\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34712\
        );

    \I__8526\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34712\
        );

    \I__8525\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34712\
        );

    \I__8524\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34712\
        );

    \I__8523\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34712\
        );

    \I__8522\ : CascadeMux
    port map (
            O => \N__34825\,
            I => \N__34708\
        );

    \I__8521\ : CascadeMux
    port map (
            O => \N__34824\,
            I => \N__34705\
        );

    \I__8520\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34686\
        );

    \I__8519\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34686\
        );

    \I__8518\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34686\
        );

    \I__8517\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34686\
        );

    \I__8516\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34686\
        );

    \I__8515\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34686\
        );

    \I__8514\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34669\
        );

    \I__8513\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34669\
        );

    \I__8512\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34669\
        );

    \I__8511\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34669\
        );

    \I__8510\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34669\
        );

    \I__8509\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34669\
        );

    \I__8508\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34669\
        );

    \I__8507\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34669\
        );

    \I__8506\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34658\
        );

    \I__8505\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34658\
        );

    \I__8504\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34658\
        );

    \I__8503\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34658\
        );

    \I__8502\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34658\
        );

    \I__8501\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34640\
        );

    \I__8500\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34640\
        );

    \I__8499\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34640\
        );

    \I__8498\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34640\
        );

    \I__8497\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34640\
        );

    \I__8496\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34640\
        );

    \I__8495\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34626\
        );

    \I__8494\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34626\
        );

    \I__8493\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34626\
        );

    \I__8492\ : CascadeMux
    port map (
            O => \N__34795\,
            I => \N__34621\
        );

    \I__8491\ : CascadeMux
    port map (
            O => \N__34794\,
            I => \N__34606\
        );

    \I__8490\ : CascadeMux
    port map (
            O => \N__34793\,
            I => \N__34603\
        );

    \I__8489\ : Span4Mux_s2_h
    port map (
            O => \N__34786\,
            I => \N__34572\
        );

    \I__8488\ : Span4Mux_s2_v
    port map (
            O => \N__34783\,
            I => \N__34572\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34572\
        );

    \I__8486\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34564\
        );

    \I__8485\ : CascadeMux
    port map (
            O => \N__34764\,
            I => \N__34561\
        );

    \I__8484\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34553\
        );

    \I__8483\ : InMux
    port map (
            O => \N__34760\,
            I => \N__34536\
        );

    \I__8482\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34536\
        );

    \I__8481\ : InMux
    port map (
            O => \N__34756\,
            I => \N__34536\
        );

    \I__8480\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34536\
        );

    \I__8479\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34536\
        );

    \I__8478\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34536\
        );

    \I__8477\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34536\
        );

    \I__8476\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34536\
        );

    \I__8475\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34521\
        );

    \I__8474\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34521\
        );

    \I__8473\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34521\
        );

    \I__8472\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34521\
        );

    \I__8471\ : InMux
    port map (
            O => \N__34744\,
            I => \N__34521\
        );

    \I__8470\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34521\
        );

    \I__8469\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34521\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__34727\,
            I => \N__34496\
        );

    \I__8467\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34491\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__34723\,
            I => \N__34488\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34485\
        );

    \I__8464\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34478\
        );

    \I__8463\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34478\
        );

    \I__8462\ : InMux
    port map (
            O => \N__34705\,
            I => \N__34478\
        );

    \I__8461\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34469\
        );

    \I__8460\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34469\
        );

    \I__8459\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34469\
        );

    \I__8458\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34469\
        );

    \I__8457\ : CascadeMux
    port map (
            O => \N__34700\,
            I => \N__34464\
        );

    \I__8456\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34461\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__34686\,
            I => \N__34454\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34454\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__34658\,
            I => \N__34454\
        );

    \I__8452\ : InMux
    port map (
            O => \N__34657\,
            I => \N__34443\
        );

    \I__8451\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34443\
        );

    \I__8450\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34443\
        );

    \I__8449\ : InMux
    port map (
            O => \N__34654\,
            I => \N__34443\
        );

    \I__8448\ : InMux
    port map (
            O => \N__34653\,
            I => \N__34443\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__34640\,
            I => \N__34440\
        );

    \I__8446\ : InMux
    port map (
            O => \N__34639\,
            I => \N__34425\
        );

    \I__8445\ : InMux
    port map (
            O => \N__34638\,
            I => \N__34425\
        );

    \I__8444\ : InMux
    port map (
            O => \N__34637\,
            I => \N__34425\
        );

    \I__8443\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34425\
        );

    \I__8442\ : InMux
    port map (
            O => \N__34635\,
            I => \N__34425\
        );

    \I__8441\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34425\
        );

    \I__8440\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34425\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__34626\,
            I => \N__34422\
        );

    \I__8438\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34409\
        );

    \I__8437\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34409\
        );

    \I__8436\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34409\
        );

    \I__8435\ : InMux
    port map (
            O => \N__34620\,
            I => \N__34409\
        );

    \I__8434\ : InMux
    port map (
            O => \N__34619\,
            I => \N__34409\
        );

    \I__8433\ : InMux
    port map (
            O => \N__34618\,
            I => \N__34409\
        );

    \I__8432\ : InMux
    port map (
            O => \N__34617\,
            I => \N__34385\
        );

    \I__8431\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34385\
        );

    \I__8430\ : InMux
    port map (
            O => \N__34615\,
            I => \N__34385\
        );

    \I__8429\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34385\
        );

    \I__8428\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34385\
        );

    \I__8427\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34385\
        );

    \I__8426\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34385\
        );

    \I__8425\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34385\
        );

    \I__8424\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34368\
        );

    \I__8423\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34368\
        );

    \I__8422\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34368\
        );

    \I__8421\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34368\
        );

    \I__8420\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34368\
        );

    \I__8419\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34368\
        );

    \I__8418\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34368\
        );

    \I__8417\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34368\
        );

    \I__8416\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34351\
        );

    \I__8415\ : InMux
    port map (
            O => \N__34596\,
            I => \N__34351\
        );

    \I__8414\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34351\
        );

    \I__8413\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34351\
        );

    \I__8412\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34351\
        );

    \I__8411\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34351\
        );

    \I__8410\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34351\
        );

    \I__8409\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34351\
        );

    \I__8408\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34334\
        );

    \I__8407\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34334\
        );

    \I__8406\ : InMux
    port map (
            O => \N__34587\,
            I => \N__34334\
        );

    \I__8405\ : InMux
    port map (
            O => \N__34586\,
            I => \N__34334\
        );

    \I__8404\ : InMux
    port map (
            O => \N__34585\,
            I => \N__34334\
        );

    \I__8403\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34334\
        );

    \I__8402\ : InMux
    port map (
            O => \N__34583\,
            I => \N__34334\
        );

    \I__8401\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34334\
        );

    \I__8400\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34327\
        );

    \I__8399\ : InMux
    port map (
            O => \N__34580\,
            I => \N__34327\
        );

    \I__8398\ : InMux
    port map (
            O => \N__34579\,
            I => \N__34327\
        );

    \I__8397\ : Span4Mux_v
    port map (
            O => \N__34572\,
            I => \N__34322\
        );

    \I__8396\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34319\
        );

    \I__8395\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34316\
        );

    \I__8394\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34313\
        );

    \I__8393\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34310\
        );

    \I__8392\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34307\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34300\
        );

    \I__8390\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34287\
        );

    \I__8389\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34287\
        );

    \I__8388\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34287\
        );

    \I__8387\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34287\
        );

    \I__8386\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34287\
        );

    \I__8385\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34287\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__34553\,
            I => \N__34280\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__34536\,
            I => \N__34280\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__34521\,
            I => \N__34280\
        );

    \I__8381\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34277\
        );

    \I__8380\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34267\
        );

    \I__8379\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34267\
        );

    \I__8378\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34267\
        );

    \I__8377\ : InMux
    port map (
            O => \N__34516\,
            I => \N__34267\
        );

    \I__8376\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34264\
        );

    \I__8375\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34247\
        );

    \I__8374\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34247\
        );

    \I__8373\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34247\
        );

    \I__8372\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34247\
        );

    \I__8371\ : InMux
    port map (
            O => \N__34510\,
            I => \N__34247\
        );

    \I__8370\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34247\
        );

    \I__8369\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34247\
        );

    \I__8368\ : InMux
    port map (
            O => \N__34507\,
            I => \N__34247\
        );

    \I__8367\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34230\
        );

    \I__8366\ : InMux
    port map (
            O => \N__34505\,
            I => \N__34230\
        );

    \I__8365\ : InMux
    port map (
            O => \N__34504\,
            I => \N__34230\
        );

    \I__8364\ : InMux
    port map (
            O => \N__34503\,
            I => \N__34230\
        );

    \I__8363\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34230\
        );

    \I__8362\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34230\
        );

    \I__8361\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34230\
        );

    \I__8360\ : InMux
    port map (
            O => \N__34499\,
            I => \N__34230\
        );

    \I__8359\ : Span4Mux_s3_h
    port map (
            O => \N__34496\,
            I => \N__34227\
        );

    \I__8358\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34222\
        );

    \I__8357\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34222\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__34491\,
            I => \N__34219\
        );

    \I__8355\ : Span4Mux_v
    port map (
            O => \N__34488\,
            I => \N__34216\
        );

    \I__8354\ : Span4Mux_v
    port map (
            O => \N__34485\,
            I => \N__34211\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__34478\,
            I => \N__34211\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__34469\,
            I => \N__34208\
        );

    \I__8351\ : CascadeMux
    port map (
            O => \N__34468\,
            I => \N__34184\
        );

    \I__8350\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34177\
        );

    \I__8349\ : InMux
    port map (
            O => \N__34464\,
            I => \N__34174\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__34461\,
            I => \N__34167\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__34454\,
            I => \N__34167\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__34443\,
            I => \N__34167\
        );

    \I__8345\ : Span4Mux_h
    port map (
            O => \N__34440\,
            I => \N__34158\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__34425\,
            I => \N__34158\
        );

    \I__8343\ : Span4Mux_s3_v
    port map (
            O => \N__34422\,
            I => \N__34158\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__34409\,
            I => \N__34158\
        );

    \I__8341\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34143\
        );

    \I__8340\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34143\
        );

    \I__8339\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34143\
        );

    \I__8338\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34143\
        );

    \I__8337\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34143\
        );

    \I__8336\ : InMux
    port map (
            O => \N__34403\,
            I => \N__34143\
        );

    \I__8335\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34143\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__34385\,
            I => \N__34134\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__34368\,
            I => \N__34134\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__34351\,
            I => \N__34134\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34134\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__34327\,
            I => \N__34131\
        );

    \I__8329\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34124\
        );

    \I__8328\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34121\
        );

    \I__8327\ : Span4Mux_h
    port map (
            O => \N__34322\,
            I => \N__34108\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__34319\,
            I => \N__34108\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__34316\,
            I => \N__34108\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__34313\,
            I => \N__34108\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__34310\,
            I => \N__34108\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__34307\,
            I => \N__34108\
        );

    \I__8321\ : InMux
    port map (
            O => \N__34306\,
            I => \N__34105\
        );

    \I__8320\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34102\
        );

    \I__8319\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34097\
        );

    \I__8318\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34097\
        );

    \I__8317\ : Span4Mux_s2_v
    port map (
            O => \N__34300\,
            I => \N__34092\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34092\
        );

    \I__8315\ : Span4Mux_v
    port map (
            O => \N__34280\,
            I => \N__34089\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34086\
        );

    \I__8313\ : CascadeMux
    port map (
            O => \N__34276\,
            I => \N__34075\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__34267\,
            I => \N__34059\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__34264\,
            I => \N__34059\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__34247\,
            I => \N__34059\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34059\
        );

    \I__8308\ : Span4Mux_v
    port map (
            O => \N__34227\,
            I => \N__34054\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__34222\,
            I => \N__34054\
        );

    \I__8306\ : Span4Mux_v
    port map (
            O => \N__34219\,
            I => \N__34045\
        );

    \I__8305\ : Span4Mux_s0_h
    port map (
            O => \N__34216\,
            I => \N__34045\
        );

    \I__8304\ : Span4Mux_v
    port map (
            O => \N__34211\,
            I => \N__34045\
        );

    \I__8303\ : Span4Mux_v
    port map (
            O => \N__34208\,
            I => \N__34045\
        );

    \I__8302\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34034\
        );

    \I__8301\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34034\
        );

    \I__8300\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34034\
        );

    \I__8299\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34034\
        );

    \I__8298\ : InMux
    port map (
            O => \N__34203\,
            I => \N__34034\
        );

    \I__8297\ : InMux
    port map (
            O => \N__34202\,
            I => \N__34023\
        );

    \I__8296\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34023\
        );

    \I__8295\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34023\
        );

    \I__8294\ : InMux
    port map (
            O => \N__34199\,
            I => \N__34023\
        );

    \I__8293\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34023\
        );

    \I__8292\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34006\
        );

    \I__8291\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34006\
        );

    \I__8290\ : InMux
    port map (
            O => \N__34195\,
            I => \N__34006\
        );

    \I__8289\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34006\
        );

    \I__8288\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34006\
        );

    \I__8287\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34006\
        );

    \I__8286\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34006\
        );

    \I__8285\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34006\
        );

    \I__8284\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34003\
        );

    \I__8283\ : InMux
    port map (
            O => \N__34188\,
            I => \N__33988\
        );

    \I__8282\ : InMux
    port map (
            O => \N__34187\,
            I => \N__33988\
        );

    \I__8281\ : InMux
    port map (
            O => \N__34184\,
            I => \N__33988\
        );

    \I__8280\ : InMux
    port map (
            O => \N__34183\,
            I => \N__33988\
        );

    \I__8279\ : InMux
    port map (
            O => \N__34182\,
            I => \N__33988\
        );

    \I__8278\ : InMux
    port map (
            O => \N__34181\,
            I => \N__33988\
        );

    \I__8277\ : InMux
    port map (
            O => \N__34180\,
            I => \N__33988\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__34177\,
            I => \N__33979\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__34174\,
            I => \N__33979\
        );

    \I__8274\ : Span4Mux_v
    port map (
            O => \N__34167\,
            I => \N__33979\
        );

    \I__8273\ : Span4Mux_v
    port map (
            O => \N__34158\,
            I => \N__33979\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__34143\,
            I => \N__33976\
        );

    \I__8271\ : Span4Mux_v
    port map (
            O => \N__34134\,
            I => \N__33971\
        );

    \I__8270\ : Span4Mux_s2_v
    port map (
            O => \N__34131\,
            I => \N__33971\
        );

    \I__8269\ : InMux
    port map (
            O => \N__34130\,
            I => \N__33968\
        );

    \I__8268\ : InMux
    port map (
            O => \N__34129\,
            I => \N__33963\
        );

    \I__8267\ : InMux
    port map (
            O => \N__34128\,
            I => \N__33963\
        );

    \I__8266\ : InMux
    port map (
            O => \N__34127\,
            I => \N__33960\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__34124\,
            I => \N__33955\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__34121\,
            I => \N__33955\
        );

    \I__8263\ : Span4Mux_s2_v
    port map (
            O => \N__34108\,
            I => \N__33932\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__34105\,
            I => \N__33932\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__34102\,
            I => \N__33932\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__34097\,
            I => \N__33932\
        );

    \I__8259\ : Span4Mux_v
    port map (
            O => \N__34092\,
            I => \N__33932\
        );

    \I__8258\ : Span4Mux_s1_h
    port map (
            O => \N__34089\,
            I => \N__33932\
        );

    \I__8257\ : Span4Mux_s2_v
    port map (
            O => \N__34086\,
            I => \N__33932\
        );

    \I__8256\ : InMux
    port map (
            O => \N__34085\,
            I => \N__33921\
        );

    \I__8255\ : InMux
    port map (
            O => \N__34084\,
            I => \N__33921\
        );

    \I__8254\ : InMux
    port map (
            O => \N__34083\,
            I => \N__33914\
        );

    \I__8253\ : InMux
    port map (
            O => \N__34082\,
            I => \N__33914\
        );

    \I__8252\ : InMux
    port map (
            O => \N__34081\,
            I => \N__33914\
        );

    \I__8251\ : InMux
    port map (
            O => \N__34080\,
            I => \N__33909\
        );

    \I__8250\ : InMux
    port map (
            O => \N__34079\,
            I => \N__33909\
        );

    \I__8249\ : CascadeMux
    port map (
            O => \N__34078\,
            I => \N__33905\
        );

    \I__8248\ : InMux
    port map (
            O => \N__34075\,
            I => \N__33899\
        );

    \I__8247\ : InMux
    port map (
            O => \N__34074\,
            I => \N__33884\
        );

    \I__8246\ : InMux
    port map (
            O => \N__34073\,
            I => \N__33884\
        );

    \I__8245\ : InMux
    port map (
            O => \N__34072\,
            I => \N__33884\
        );

    \I__8244\ : InMux
    port map (
            O => \N__34071\,
            I => \N__33884\
        );

    \I__8243\ : InMux
    port map (
            O => \N__34070\,
            I => \N__33884\
        );

    \I__8242\ : InMux
    port map (
            O => \N__34069\,
            I => \N__33884\
        );

    \I__8241\ : InMux
    port map (
            O => \N__34068\,
            I => \N__33884\
        );

    \I__8240\ : Span4Mux_v
    port map (
            O => \N__34059\,
            I => \N__33879\
        );

    \I__8239\ : Span4Mux_h
    port map (
            O => \N__34054\,
            I => \N__33879\
        );

    \I__8238\ : Sp12to4
    port map (
            O => \N__34045\,
            I => \N__33870\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__34034\,
            I => \N__33870\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__34023\,
            I => \N__33870\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__34006\,
            I => \N__33870\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__34003\,
            I => \N__33866\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__33988\,
            I => \N__33863\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__33979\,
            I => \N__33858\
        );

    \I__8231\ : Span4Mux_h
    port map (
            O => \N__33976\,
            I => \N__33858\
        );

    \I__8230\ : Sp12to4
    port map (
            O => \N__33971\,
            I => \N__33855\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__33968\,
            I => \N__33846\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__33963\,
            I => \N__33846\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__33960\,
            I => \N__33846\
        );

    \I__8226\ : Span4Mux_h
    port map (
            O => \N__33955\,
            I => \N__33846\
        );

    \I__8225\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33829\
        );

    \I__8224\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33829\
        );

    \I__8223\ : InMux
    port map (
            O => \N__33952\,
            I => \N__33829\
        );

    \I__8222\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33829\
        );

    \I__8221\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33829\
        );

    \I__8220\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33829\
        );

    \I__8219\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33829\
        );

    \I__8218\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33829\
        );

    \I__8217\ : Sp12to4
    port map (
            O => \N__33932\,
            I => \N__33826\
        );

    \I__8216\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33810\
        );

    \I__8215\ : InMux
    port map (
            O => \N__33930\,
            I => \N__33810\
        );

    \I__8214\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33810\
        );

    \I__8213\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33810\
        );

    \I__8212\ : InMux
    port map (
            O => \N__33927\,
            I => \N__33810\
        );

    \I__8211\ : InMux
    port map (
            O => \N__33926\,
            I => \N__33810\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__33921\,
            I => \N__33803\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__33914\,
            I => \N__33803\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__33909\,
            I => \N__33803\
        );

    \I__8207\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33792\
        );

    \I__8206\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33792\
        );

    \I__8205\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33792\
        );

    \I__8204\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33792\
        );

    \I__8203\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33792\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33787\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__33884\,
            I => \N__33787\
        );

    \I__8200\ : Sp12to4
    port map (
            O => \N__33879\,
            I => \N__33782\
        );

    \I__8199\ : Span12Mux_s7_h
    port map (
            O => \N__33870\,
            I => \N__33782\
        );

    \I__8198\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33779\
        );

    \I__8197\ : Span4Mux_h
    port map (
            O => \N__33866\,
            I => \N__33772\
        );

    \I__8196\ : Span4Mux_h
    port map (
            O => \N__33863\,
            I => \N__33772\
        );

    \I__8195\ : Span4Mux_v
    port map (
            O => \N__33858\,
            I => \N__33772\
        );

    \I__8194\ : Span12Mux_s7_h
    port map (
            O => \N__33855\,
            I => \N__33763\
        );

    \I__8193\ : Sp12to4
    port map (
            O => \N__33846\,
            I => \N__33763\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__33829\,
            I => \N__33763\
        );

    \I__8191\ : Span12Mux_s4_h
    port map (
            O => \N__33826\,
            I => \N__33763\
        );

    \I__8190\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33760\
        );

    \I__8189\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33755\
        );

    \I__8188\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33755\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__33810\,
            I => \N__33750\
        );

    \I__8186\ : Span12Mux_v
    port map (
            O => \N__33803\,
            I => \N__33750\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__33792\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__33787\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8183\ : Odrv12
    port map (
            O => \N__33782\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__33779\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8181\ : Odrv4
    port map (
            O => \N__33772\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8180\ : Odrv12
    port map (
            O => \N__33763\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__33760\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__33755\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8177\ : Odrv12
    port map (
            O => \N__33750\,
            I => \processor_zipi8.alu_mux_sel_0\
        );

    \I__8176\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33727\
        );

    \I__8175\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33724\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__33727\,
            I => \N__33719\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__33724\,
            I => \N__33719\
        );

    \I__8172\ : Span4Mux_h
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__8171\ : Span4Mux_h
    port map (
            O => \N__33716\,
            I => \N__33713\
        );

    \I__8170\ : Odrv4
    port map (
            O => \N__33713\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_4\
        );

    \I__8169\ : ClkMux
    port map (
            O => \N__33710\,
            I => \N__33395\
        );

    \I__8168\ : ClkMux
    port map (
            O => \N__33709\,
            I => \N__33395\
        );

    \I__8167\ : ClkMux
    port map (
            O => \N__33708\,
            I => \N__33395\
        );

    \I__8166\ : ClkMux
    port map (
            O => \N__33707\,
            I => \N__33395\
        );

    \I__8165\ : ClkMux
    port map (
            O => \N__33706\,
            I => \N__33395\
        );

    \I__8164\ : ClkMux
    port map (
            O => \N__33705\,
            I => \N__33395\
        );

    \I__8163\ : ClkMux
    port map (
            O => \N__33704\,
            I => \N__33395\
        );

    \I__8162\ : ClkMux
    port map (
            O => \N__33703\,
            I => \N__33395\
        );

    \I__8161\ : ClkMux
    port map (
            O => \N__33702\,
            I => \N__33395\
        );

    \I__8160\ : ClkMux
    port map (
            O => \N__33701\,
            I => \N__33395\
        );

    \I__8159\ : ClkMux
    port map (
            O => \N__33700\,
            I => \N__33395\
        );

    \I__8158\ : ClkMux
    port map (
            O => \N__33699\,
            I => \N__33395\
        );

    \I__8157\ : ClkMux
    port map (
            O => \N__33698\,
            I => \N__33395\
        );

    \I__8156\ : ClkMux
    port map (
            O => \N__33697\,
            I => \N__33395\
        );

    \I__8155\ : ClkMux
    port map (
            O => \N__33696\,
            I => \N__33395\
        );

    \I__8154\ : ClkMux
    port map (
            O => \N__33695\,
            I => \N__33395\
        );

    \I__8153\ : ClkMux
    port map (
            O => \N__33694\,
            I => \N__33395\
        );

    \I__8152\ : ClkMux
    port map (
            O => \N__33693\,
            I => \N__33395\
        );

    \I__8151\ : ClkMux
    port map (
            O => \N__33692\,
            I => \N__33395\
        );

    \I__8150\ : ClkMux
    port map (
            O => \N__33691\,
            I => \N__33395\
        );

    \I__8149\ : ClkMux
    port map (
            O => \N__33690\,
            I => \N__33395\
        );

    \I__8148\ : ClkMux
    port map (
            O => \N__33689\,
            I => \N__33395\
        );

    \I__8147\ : ClkMux
    port map (
            O => \N__33688\,
            I => \N__33395\
        );

    \I__8146\ : ClkMux
    port map (
            O => \N__33687\,
            I => \N__33395\
        );

    \I__8145\ : ClkMux
    port map (
            O => \N__33686\,
            I => \N__33395\
        );

    \I__8144\ : ClkMux
    port map (
            O => \N__33685\,
            I => \N__33395\
        );

    \I__8143\ : ClkMux
    port map (
            O => \N__33684\,
            I => \N__33395\
        );

    \I__8142\ : ClkMux
    port map (
            O => \N__33683\,
            I => \N__33395\
        );

    \I__8141\ : ClkMux
    port map (
            O => \N__33682\,
            I => \N__33395\
        );

    \I__8140\ : ClkMux
    port map (
            O => \N__33681\,
            I => \N__33395\
        );

    \I__8139\ : ClkMux
    port map (
            O => \N__33680\,
            I => \N__33395\
        );

    \I__8138\ : ClkMux
    port map (
            O => \N__33679\,
            I => \N__33395\
        );

    \I__8137\ : ClkMux
    port map (
            O => \N__33678\,
            I => \N__33395\
        );

    \I__8136\ : ClkMux
    port map (
            O => \N__33677\,
            I => \N__33395\
        );

    \I__8135\ : ClkMux
    port map (
            O => \N__33676\,
            I => \N__33395\
        );

    \I__8134\ : ClkMux
    port map (
            O => \N__33675\,
            I => \N__33395\
        );

    \I__8133\ : ClkMux
    port map (
            O => \N__33674\,
            I => \N__33395\
        );

    \I__8132\ : ClkMux
    port map (
            O => \N__33673\,
            I => \N__33395\
        );

    \I__8131\ : ClkMux
    port map (
            O => \N__33672\,
            I => \N__33395\
        );

    \I__8130\ : ClkMux
    port map (
            O => \N__33671\,
            I => \N__33395\
        );

    \I__8129\ : ClkMux
    port map (
            O => \N__33670\,
            I => \N__33395\
        );

    \I__8128\ : ClkMux
    port map (
            O => \N__33669\,
            I => \N__33395\
        );

    \I__8127\ : ClkMux
    port map (
            O => \N__33668\,
            I => \N__33395\
        );

    \I__8126\ : ClkMux
    port map (
            O => \N__33667\,
            I => \N__33395\
        );

    \I__8125\ : ClkMux
    port map (
            O => \N__33666\,
            I => \N__33395\
        );

    \I__8124\ : ClkMux
    port map (
            O => \N__33665\,
            I => \N__33395\
        );

    \I__8123\ : ClkMux
    port map (
            O => \N__33664\,
            I => \N__33395\
        );

    \I__8122\ : ClkMux
    port map (
            O => \N__33663\,
            I => \N__33395\
        );

    \I__8121\ : ClkMux
    port map (
            O => \N__33662\,
            I => \N__33395\
        );

    \I__8120\ : ClkMux
    port map (
            O => \N__33661\,
            I => \N__33395\
        );

    \I__8119\ : ClkMux
    port map (
            O => \N__33660\,
            I => \N__33395\
        );

    \I__8118\ : ClkMux
    port map (
            O => \N__33659\,
            I => \N__33395\
        );

    \I__8117\ : ClkMux
    port map (
            O => \N__33658\,
            I => \N__33395\
        );

    \I__8116\ : ClkMux
    port map (
            O => \N__33657\,
            I => \N__33395\
        );

    \I__8115\ : ClkMux
    port map (
            O => \N__33656\,
            I => \N__33395\
        );

    \I__8114\ : ClkMux
    port map (
            O => \N__33655\,
            I => \N__33395\
        );

    \I__8113\ : ClkMux
    port map (
            O => \N__33654\,
            I => \N__33395\
        );

    \I__8112\ : ClkMux
    port map (
            O => \N__33653\,
            I => \N__33395\
        );

    \I__8111\ : ClkMux
    port map (
            O => \N__33652\,
            I => \N__33395\
        );

    \I__8110\ : ClkMux
    port map (
            O => \N__33651\,
            I => \N__33395\
        );

    \I__8109\ : ClkMux
    port map (
            O => \N__33650\,
            I => \N__33395\
        );

    \I__8108\ : ClkMux
    port map (
            O => \N__33649\,
            I => \N__33395\
        );

    \I__8107\ : ClkMux
    port map (
            O => \N__33648\,
            I => \N__33395\
        );

    \I__8106\ : ClkMux
    port map (
            O => \N__33647\,
            I => \N__33395\
        );

    \I__8105\ : ClkMux
    port map (
            O => \N__33646\,
            I => \N__33395\
        );

    \I__8104\ : ClkMux
    port map (
            O => \N__33645\,
            I => \N__33395\
        );

    \I__8103\ : ClkMux
    port map (
            O => \N__33644\,
            I => \N__33395\
        );

    \I__8102\ : ClkMux
    port map (
            O => \N__33643\,
            I => \N__33395\
        );

    \I__8101\ : ClkMux
    port map (
            O => \N__33642\,
            I => \N__33395\
        );

    \I__8100\ : ClkMux
    port map (
            O => \N__33641\,
            I => \N__33395\
        );

    \I__8099\ : ClkMux
    port map (
            O => \N__33640\,
            I => \N__33395\
        );

    \I__8098\ : ClkMux
    port map (
            O => \N__33639\,
            I => \N__33395\
        );

    \I__8097\ : ClkMux
    port map (
            O => \N__33638\,
            I => \N__33395\
        );

    \I__8096\ : ClkMux
    port map (
            O => \N__33637\,
            I => \N__33395\
        );

    \I__8095\ : ClkMux
    port map (
            O => \N__33636\,
            I => \N__33395\
        );

    \I__8094\ : ClkMux
    port map (
            O => \N__33635\,
            I => \N__33395\
        );

    \I__8093\ : ClkMux
    port map (
            O => \N__33634\,
            I => \N__33395\
        );

    \I__8092\ : ClkMux
    port map (
            O => \N__33633\,
            I => \N__33395\
        );

    \I__8091\ : ClkMux
    port map (
            O => \N__33632\,
            I => \N__33395\
        );

    \I__8090\ : ClkMux
    port map (
            O => \N__33631\,
            I => \N__33395\
        );

    \I__8089\ : ClkMux
    port map (
            O => \N__33630\,
            I => \N__33395\
        );

    \I__8088\ : ClkMux
    port map (
            O => \N__33629\,
            I => \N__33395\
        );

    \I__8087\ : ClkMux
    port map (
            O => \N__33628\,
            I => \N__33395\
        );

    \I__8086\ : ClkMux
    port map (
            O => \N__33627\,
            I => \N__33395\
        );

    \I__8085\ : ClkMux
    port map (
            O => \N__33626\,
            I => \N__33395\
        );

    \I__8084\ : ClkMux
    port map (
            O => \N__33625\,
            I => \N__33395\
        );

    \I__8083\ : ClkMux
    port map (
            O => \N__33624\,
            I => \N__33395\
        );

    \I__8082\ : ClkMux
    port map (
            O => \N__33623\,
            I => \N__33395\
        );

    \I__8081\ : ClkMux
    port map (
            O => \N__33622\,
            I => \N__33395\
        );

    \I__8080\ : ClkMux
    port map (
            O => \N__33621\,
            I => \N__33395\
        );

    \I__8079\ : ClkMux
    port map (
            O => \N__33620\,
            I => \N__33395\
        );

    \I__8078\ : ClkMux
    port map (
            O => \N__33619\,
            I => \N__33395\
        );

    \I__8077\ : ClkMux
    port map (
            O => \N__33618\,
            I => \N__33395\
        );

    \I__8076\ : ClkMux
    port map (
            O => \N__33617\,
            I => \N__33395\
        );

    \I__8075\ : ClkMux
    port map (
            O => \N__33616\,
            I => \N__33395\
        );

    \I__8074\ : ClkMux
    port map (
            O => \N__33615\,
            I => \N__33395\
        );

    \I__8073\ : ClkMux
    port map (
            O => \N__33614\,
            I => \N__33395\
        );

    \I__8072\ : ClkMux
    port map (
            O => \N__33613\,
            I => \N__33395\
        );

    \I__8071\ : ClkMux
    port map (
            O => \N__33612\,
            I => \N__33395\
        );

    \I__8070\ : ClkMux
    port map (
            O => \N__33611\,
            I => \N__33395\
        );

    \I__8069\ : ClkMux
    port map (
            O => \N__33610\,
            I => \N__33395\
        );

    \I__8068\ : ClkMux
    port map (
            O => \N__33609\,
            I => \N__33395\
        );

    \I__8067\ : ClkMux
    port map (
            O => \N__33608\,
            I => \N__33395\
        );

    \I__8066\ : ClkMux
    port map (
            O => \N__33607\,
            I => \N__33395\
        );

    \I__8065\ : ClkMux
    port map (
            O => \N__33606\,
            I => \N__33395\
        );

    \I__8064\ : GlobalMux
    port map (
            O => \N__33395\,
            I => \N__33392\
        );

    \I__8063\ : gio2CtrlBuf
    port map (
            O => \N__33392\,
            I => \CLK_3P3_MHZ_c_g\
        );

    \I__8062\ : CEMux
    port map (
            O => \N__33389\,
            I => \N__33386\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__33386\,
            I => \N__33382\
        );

    \I__8060\ : CEMux
    port map (
            O => \N__33385\,
            I => \N__33379\
        );

    \I__8059\ : Span4Mux_s0_h
    port map (
            O => \N__33382\,
            I => \N__33376\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__33379\,
            I => \N__33373\
        );

    \I__8057\ : Span4Mux_h
    port map (
            O => \N__33376\,
            I => \N__33370\
        );

    \I__8056\ : Span4Mux_s3_v
    port map (
            O => \N__33373\,
            I => \N__33367\
        );

    \I__8055\ : Span4Mux_v
    port map (
            O => \N__33370\,
            I => \N__33364\
        );

    \I__8054\ : Odrv4
    port map (
            O => \N__33367\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22\
        );

    \I__8053\ : Odrv4
    port map (
            O => \N__33364\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22\
        );

    \I__8052\ : CascadeMux
    port map (
            O => \N__33359\,
            I => \N__33355\
        );

    \I__8051\ : InMux
    port map (
            O => \N__33358\,
            I => \N__33352\
        );

    \I__8050\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33349\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__33352\,
            I => \N__33346\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__33349\,
            I => \N__33343\
        );

    \I__8047\ : Span4Mux_h
    port map (
            O => \N__33346\,
            I => \N__33328\
        );

    \I__8046\ : Span4Mux_s3_h
    port map (
            O => \N__33343\,
            I => \N__33328\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__33342\,
            I => \N__33324\
        );

    \I__8044\ : CascadeMux
    port map (
            O => \N__33341\,
            I => \N__33321\
        );

    \I__8043\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33313\
        );

    \I__8042\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33306\
        );

    \I__8041\ : InMux
    port map (
            O => \N__33338\,
            I => \N__33303\
        );

    \I__8040\ : CascadeMux
    port map (
            O => \N__33337\,
            I => \N__33298\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__33336\,
            I => \N__33295\
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__33335\,
            I => \N__33291\
        );

    \I__8037\ : InMux
    port map (
            O => \N__33334\,
            I => \N__33287\
        );

    \I__8036\ : InMux
    port map (
            O => \N__33333\,
            I => \N__33284\
        );

    \I__8035\ : IoSpan4Mux
    port map (
            O => \N__33328\,
            I => \N__33281\
        );

    \I__8034\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33278\
        );

    \I__8033\ : InMux
    port map (
            O => \N__33324\,
            I => \N__33275\
        );

    \I__8032\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33272\
        );

    \I__8031\ : CascadeMux
    port map (
            O => \N__33320\,
            I => \N__33267\
        );

    \I__8030\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33263\
        );

    \I__8029\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33260\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__33317\,
            I => \N__33257\
        );

    \I__8027\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33253\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33250\
        );

    \I__8025\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33247\
        );

    \I__8024\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33244\
        );

    \I__8023\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33241\
        );

    \I__8022\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33238\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__33306\,
            I => \N__33235\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__33303\,
            I => \N__33232\
        );

    \I__8019\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33229\
        );

    \I__8018\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33226\
        );

    \I__8017\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33223\
        );

    \I__8016\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33220\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__33294\,
            I => \N__33216\
        );

    \I__8014\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33213\
        );

    \I__8013\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33210\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__33287\,
            I => \N__33207\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__33284\,
            I => \N__33204\
        );

    \I__8010\ : Span4Mux_s0_v
    port map (
            O => \N__33281\,
            I => \N__33194\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33194\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__33275\,
            I => \N__33194\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__33272\,
            I => \N__33194\
        );

    \I__8006\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33191\
        );

    \I__8005\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33186\
        );

    \I__8004\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33186\
        );

    \I__8003\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33183\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__33263\,
            I => \N__33178\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__33260\,
            I => \N__33178\
        );

    \I__8000\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33175\
        );

    \I__7999\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33171\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__33253\,
            I => \N__33164\
        );

    \I__7997\ : Span4Mux_v
    port map (
            O => \N__33250\,
            I => \N__33164\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__33247\,
            I => \N__33164\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__33244\,
            I => \N__33161\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33148\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33148\
        );

    \I__7992\ : Span4Mux_s3_h
    port map (
            O => \N__33235\,
            I => \N__33148\
        );

    \I__7991\ : Span4Mux_v
    port map (
            O => \N__33232\,
            I => \N__33148\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__33229\,
            I => \N__33148\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__33226\,
            I => \N__33148\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__33223\,
            I => \N__33142\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__33220\,
            I => \N__33142\
        );

    \I__7986\ : InMux
    port map (
            O => \N__33219\,
            I => \N__33139\
        );

    \I__7985\ : InMux
    port map (
            O => \N__33216\,
            I => \N__33136\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__33213\,
            I => \N__33133\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__33210\,
            I => \N__33130\
        );

    \I__7982\ : Span4Mux_v
    port map (
            O => \N__33207\,
            I => \N__33125\
        );

    \I__7981\ : Span4Mux_s0_h
    port map (
            O => \N__33204\,
            I => \N__33125\
        );

    \I__7980\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33122\
        );

    \I__7979\ : Span4Mux_h
    port map (
            O => \N__33194\,
            I => \N__33119\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33114\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__33186\,
            I => \N__33114\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33111\
        );

    \I__7975\ : Span4Mux_v
    port map (
            O => \N__33178\,
            I => \N__33108\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__33175\,
            I => \N__33105\
        );

    \I__7973\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33102\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__33171\,
            I => \N__33093\
        );

    \I__7971\ : Span4Mux_h
    port map (
            O => \N__33164\,
            I => \N__33093\
        );

    \I__7970\ : Span4Mux_s1_v
    port map (
            O => \N__33161\,
            I => \N__33093\
        );

    \I__7969\ : Span4Mux_h
    port map (
            O => \N__33148\,
            I => \N__33093\
        );

    \I__7968\ : CascadeMux
    port map (
            O => \N__33147\,
            I => \N__33090\
        );

    \I__7967\ : Span4Mux_v
    port map (
            O => \N__33142\,
            I => \N__33087\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__33139\,
            I => \N__33080\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__33136\,
            I => \N__33080\
        );

    \I__7964\ : Span4Mux_s3_v
    port map (
            O => \N__33133\,
            I => \N__33080\
        );

    \I__7963\ : Span4Mux_v
    port map (
            O => \N__33130\,
            I => \N__33077\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__33125\,
            I => \N__33072\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__33122\,
            I => \N__33072\
        );

    \I__7960\ : Span4Mux_v
    port map (
            O => \N__33119\,
            I => \N__33067\
        );

    \I__7959\ : Span4Mux_s3_h
    port map (
            O => \N__33114\,
            I => \N__33067\
        );

    \I__7958\ : Span4Mux_v
    port map (
            O => \N__33111\,
            I => \N__33062\
        );

    \I__7957\ : Span4Mux_s1_h
    port map (
            O => \N__33108\,
            I => \N__33062\
        );

    \I__7956\ : Span12Mux_s7_h
    port map (
            O => \N__33105\,
            I => \N__33059\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__33102\,
            I => \N__33054\
        );

    \I__7954\ : Span4Mux_v
    port map (
            O => \N__33093\,
            I => \N__33054\
        );

    \I__7953\ : InMux
    port map (
            O => \N__33090\,
            I => \N__33051\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__33087\,
            I => \N__33040\
        );

    \I__7951\ : Span4Mux_v
    port map (
            O => \N__33080\,
            I => \N__33040\
        );

    \I__7950\ : Span4Mux_h
    port map (
            O => \N__33077\,
            I => \N__33040\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__33072\,
            I => \N__33040\
        );

    \I__7948\ : Span4Mux_v
    port map (
            O => \N__33067\,
            I => \N__33040\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__33062\,
            I => \processor_zipi8.arith_logical_result_7\
        );

    \I__7946\ : Odrv12
    port map (
            O => \N__33059\,
            I => \processor_zipi8.arith_logical_result_7\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__33054\,
            I => \processor_zipi8.arith_logical_result_7\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__33051\,
            I => \processor_zipi8.arith_logical_result_7\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__33040\,
            I => \processor_zipi8.arith_logical_result_7\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__33029\,
            I => \N__33025\
        );

    \I__7941\ : CascadeMux
    port map (
            O => \N__33028\,
            I => \N__33022\
        );

    \I__7940\ : InMux
    port map (
            O => \N__33025\,
            I => \N__33018\
        );

    \I__7939\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33006\
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__33021\,
            I => \N__33003\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__33018\,
            I => \N__32996\
        );

    \I__7936\ : CascadeMux
    port map (
            O => \N__33017\,
            I => \N__32990\
        );

    \I__7935\ : InMux
    port map (
            O => \N__33016\,
            I => \N__32987\
        );

    \I__7934\ : InMux
    port map (
            O => \N__33015\,
            I => \N__32984\
        );

    \I__7933\ : CascadeMux
    port map (
            O => \N__33014\,
            I => \N__32981\
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__33013\,
            I => \N__32975\
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__33012\,
            I => \N__32970\
        );

    \I__7930\ : CascadeMux
    port map (
            O => \N__33011\,
            I => \N__32967\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__33010\,
            I => \N__32964\
        );

    \I__7928\ : CascadeMux
    port map (
            O => \N__33009\,
            I => \N__32961\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__33006\,
            I => \N__32957\
        );

    \I__7926\ : InMux
    port map (
            O => \N__33003\,
            I => \N__32954\
        );

    \I__7925\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32951\
        );

    \I__7924\ : CascadeMux
    port map (
            O => \N__33001\,
            I => \N__32948\
        );

    \I__7923\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32945\
        );

    \I__7922\ : CascadeMux
    port map (
            O => \N__32999\,
            I => \N__32941\
        );

    \I__7921\ : Span4Mux_v
    port map (
            O => \N__32996\,
            I => \N__32938\
        );

    \I__7920\ : CascadeMux
    port map (
            O => \N__32995\,
            I => \N__32935\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__32994\,
            I => \N__32932\
        );

    \I__7918\ : InMux
    port map (
            O => \N__32993\,
            I => \N__32929\
        );

    \I__7917\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32926\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__32987\,
            I => \N__32923\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__32984\,
            I => \N__32920\
        );

    \I__7914\ : InMux
    port map (
            O => \N__32981\,
            I => \N__32917\
        );

    \I__7913\ : InMux
    port map (
            O => \N__32980\,
            I => \N__32914\
        );

    \I__7912\ : InMux
    port map (
            O => \N__32979\,
            I => \N__32911\
        );

    \I__7911\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32908\
        );

    \I__7910\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32905\
        );

    \I__7909\ : InMux
    port map (
            O => \N__32974\,
            I => \N__32902\
        );

    \I__7908\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32899\
        );

    \I__7907\ : InMux
    port map (
            O => \N__32970\,
            I => \N__32895\
        );

    \I__7906\ : InMux
    port map (
            O => \N__32967\,
            I => \N__32892\
        );

    \I__7905\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32889\
        );

    \I__7904\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32886\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__32960\,
            I => \N__32883\
        );

    \I__7902\ : Span4Mux_h
    port map (
            O => \N__32957\,
            I => \N__32876\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__32954\,
            I => \N__32876\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__32951\,
            I => \N__32876\
        );

    \I__7899\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32873\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32869\
        );

    \I__7897\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32866\
        );

    \I__7896\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32863\
        );

    \I__7895\ : Span4Mux_v
    port map (
            O => \N__32938\,
            I => \N__32860\
        );

    \I__7894\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32857\
        );

    \I__7893\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32854\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__32929\,
            I => \N__32849\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__32926\,
            I => \N__32849\
        );

    \I__7890\ : Span4Mux_s0_v
    port map (
            O => \N__32923\,
            I => \N__32838\
        );

    \I__7889\ : Span4Mux_s0_v
    port map (
            O => \N__32920\,
            I => \N__32838\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__32917\,
            I => \N__32838\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32838\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__32911\,
            I => \N__32838\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__32908\,
            I => \N__32835\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32828\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__32902\,
            I => \N__32828\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__32899\,
            I => \N__32828\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__32898\,
            I => \N__32825\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32820\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__32892\,
            I => \N__32817\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__32889\,
            I => \N__32812\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32812\
        );

    \I__7876\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32809\
        );

    \I__7875\ : Span4Mux_s3_v
    port map (
            O => \N__32876\,
            I => \N__32804\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__32873\,
            I => \N__32804\
        );

    \I__7873\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32801\
        );

    \I__7872\ : Span4Mux_s0_h
    port map (
            O => \N__32869\,
            I => \N__32794\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__32866\,
            I => \N__32794\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__32863\,
            I => \N__32794\
        );

    \I__7869\ : Span4Mux_h
    port map (
            O => \N__32860\,
            I => \N__32777\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32777\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__32854\,
            I => \N__32777\
        );

    \I__7866\ : Span4Mux_v
    port map (
            O => \N__32849\,
            I => \N__32777\
        );

    \I__7865\ : Span4Mux_v
    port map (
            O => \N__32838\,
            I => \N__32777\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__32835\,
            I => \N__32777\
        );

    \I__7863\ : Span4Mux_v
    port map (
            O => \N__32828\,
            I => \N__32777\
        );

    \I__7862\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32772\
        );

    \I__7861\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32772\
        );

    \I__7860\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32769\
        );

    \I__7859\ : Span4Mux_h
    port map (
            O => \N__32820\,
            I => \N__32762\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__32817\,
            I => \N__32762\
        );

    \I__7857\ : Span4Mux_h
    port map (
            O => \N__32812\,
            I => \N__32762\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__32809\,
            I => \N__32755\
        );

    \I__7855\ : Span4Mux_h
    port map (
            O => \N__32804\,
            I => \N__32755\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32755\
        );

    \I__7853\ : Span4Mux_v
    port map (
            O => \N__32794\,
            I => \N__32752\
        );

    \I__7852\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32749\
        );

    \I__7851\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32746\
        );

    \I__7850\ : Sp12to4
    port map (
            O => \N__32777\,
            I => \N__32741\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32741\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__32769\,
            I => \N__32736\
        );

    \I__7847\ : Span4Mux_v
    port map (
            O => \N__32762\,
            I => \N__32736\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__32755\,
            I => \N__32733\
        );

    \I__7845\ : Span4Mux_h
    port map (
            O => \N__32752\,
            I => \N__32730\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__32749\,
            I => \N__32723\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__32746\,
            I => \N__32723\
        );

    \I__7842\ : Span12Mux_s7_h
    port map (
            O => \N__32741\,
            I => \N__32723\
        );

    \I__7841\ : Odrv4
    port map (
            O => \N__32736\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__32733\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269\
        );

    \I__7839\ : Odrv4
    port map (
            O => \N__32730\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269\
        );

    \I__7838\ : Odrv12
    port map (
            O => \N__32723\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__32714\,
            I => \N__32711\
        );

    \I__7836\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32708\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32705\
        );

    \I__7834\ : Span4Mux_s2_v
    port map (
            O => \N__32705\,
            I => \N__32702\
        );

    \I__7833\ : Span4Mux_v
    port map (
            O => \N__32702\,
            I => \N__32698\
        );

    \I__7832\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32695\
        );

    \I__7831\ : Span4Mux_h
    port map (
            O => \N__32698\,
            I => \N__32692\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__32695\,
            I => \N__32689\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__32692\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7\
        );

    \I__7828\ : Odrv12
    port map (
            O => \N__32689\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7\
        );

    \I__7827\ : CEMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32678\
        );

    \I__7825\ : Span4Mux_v
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__7824\ : IoSpan4Mux
    port map (
            O => \N__32675\,
            I => \N__32671\
        );

    \I__7823\ : CEMux
    port map (
            O => \N__32674\,
            I => \N__32668\
        );

    \I__7822\ : IoSpan4Mux
    port map (
            O => \N__32671\,
            I => \N__32665\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__32668\,
            I => \N__32662\
        );

    \I__7820\ : Span4Mux_s2_h
    port map (
            O => \N__32665\,
            I => \N__32659\
        );

    \I__7819\ : Span12Mux_s3_v
    port map (
            O => \N__32662\,
            I => \N__32656\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__32659\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21\
        );

    \I__7817\ : Odrv12
    port map (
            O => \N__32656\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21\
        );

    \I__7816\ : CascadeMux
    port map (
            O => \N__32651\,
            I => \N__32647\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__32650\,
            I => \N__32644\
        );

    \I__7814\ : InMux
    port map (
            O => \N__32647\,
            I => \N__32641\
        );

    \I__7813\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32638\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32635\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32632\
        );

    \I__7810\ : Span4Mux_h
    port map (
            O => \N__32635\,
            I => \N__32629\
        );

    \I__7809\ : Span12Mux_s9_v
    port map (
            O => \N__32632\,
            I => \N__32626\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__32629\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0\
        );

    \I__7807\ : Odrv12
    port map (
            O => \N__32626\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0\
        );

    \I__7806\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32617\
        );

    \I__7805\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32614\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__32617\,
            I => \N__32611\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__32614\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1\
        );

    \I__7802\ : Odrv4
    port map (
            O => \N__32611\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1\
        );

    \I__7801\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32602\
        );

    \I__7800\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32599\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__32602\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__32599\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1\
        );

    \I__7797\ : InMux
    port map (
            O => \N__32594\,
            I => \N__32591\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__32591\,
            I => \N__32588\
        );

    \I__7795\ : Odrv12
    port map (
            O => \N__32588\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_1\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__32585\,
            I => \N__32582\
        );

    \I__7793\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32578\
        );

    \I__7792\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32575\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__32578\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__32575\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2\
        );

    \I__7789\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32566\
        );

    \I__7788\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32563\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__32566\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__32563\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2\
        );

    \I__7785\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32555\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__32555\,
            I => \N__32552\
        );

    \I__7783\ : Span4Mux_h
    port map (
            O => \N__32552\,
            I => \N__32549\
        );

    \I__7782\ : Odrv4
    port map (
            O => \N__32549\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_2\
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__32546\,
            I => \N__32542\
        );

    \I__7780\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32539\
        );

    \I__7779\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32536\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32531\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__32536\,
            I => \N__32531\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__32531\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_3\
        );

    \I__7775\ : CascadeMux
    port map (
            O => \N__32528\,
            I => \N__32525\
        );

    \I__7774\ : InMux
    port map (
            O => \N__32525\,
            I => \N__32519\
        );

    \I__7773\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32519\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__32519\,
            I => \N__32516\
        );

    \I__7771\ : Span4Mux_v
    port map (
            O => \N__32516\,
            I => \N__32513\
        );

    \I__7770\ : Span4Mux_h
    port map (
            O => \N__32513\,
            I => \N__32510\
        );

    \I__7769\ : Odrv4
    port map (
            O => \N__32510\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_4\
        );

    \I__7768\ : CEMux
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32501\
        );

    \I__7766\ : Span4Mux_s2_h
    port map (
            O => \N__32501\,
            I => \N__32498\
        );

    \I__7765\ : Span4Mux_h
    port map (
            O => \N__32498\,
            I => \N__32494\
        );

    \I__7764\ : CEMux
    port map (
            O => \N__32497\,
            I => \N__32491\
        );

    \I__7763\ : Span4Mux_v
    port map (
            O => \N__32494\,
            I => \N__32488\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32485\
        );

    \I__7761\ : Sp12to4
    port map (
            O => \N__32488\,
            I => \N__32482\
        );

    \I__7760\ : Odrv4
    port map (
            O => \N__32485\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20\
        );

    \I__7759\ : Odrv12
    port map (
            O => \N__32482\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20\
        );

    \I__7758\ : CascadeMux
    port map (
            O => \N__32477\,
            I => \N__32471\
        );

    \I__7757\ : CascadeMux
    port map (
            O => \N__32476\,
            I => \N__32468\
        );

    \I__7756\ : CascadeMux
    port map (
            O => \N__32475\,
            I => \N__32465\
        );

    \I__7755\ : CascadeMux
    port map (
            O => \N__32474\,
            I => \N__32462\
        );

    \I__7754\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32455\
        );

    \I__7753\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32452\
        );

    \I__7752\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32449\
        );

    \I__7751\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32446\
        );

    \I__7750\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32443\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__32460\,
            I => \N__32440\
        );

    \I__7748\ : CascadeMux
    port map (
            O => \N__32459\,
            I => \N__32434\
        );

    \I__7747\ : CascadeMux
    port map (
            O => \N__32458\,
            I => \N__32428\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__32455\,
            I => \N__32423\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__32452\,
            I => \N__32423\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__32449\,
            I => \N__32416\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__32446\,
            I => \N__32416\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__32443\,
            I => \N__32416\
        );

    \I__7741\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32413\
        );

    \I__7740\ : CascadeMux
    port map (
            O => \N__32439\,
            I => \N__32410\
        );

    \I__7739\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32407\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__32437\,
            I => \N__32404\
        );

    \I__7737\ : InMux
    port map (
            O => \N__32434\,
            I => \N__32400\
        );

    \I__7736\ : CascadeMux
    port map (
            O => \N__32433\,
            I => \N__32395\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__32432\,
            I => \N__32392\
        );

    \I__7734\ : CascadeMux
    port map (
            O => \N__32431\,
            I => \N__32389\
        );

    \I__7733\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32386\
        );

    \I__7732\ : Span4Mux_v
    port map (
            O => \N__32423\,
            I => \N__32381\
        );

    \I__7731\ : Span4Mux_v
    port map (
            O => \N__32416\,
            I => \N__32381\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__32413\,
            I => \N__32377\
        );

    \I__7729\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32374\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32371\
        );

    \I__7727\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32368\
        );

    \I__7726\ : CascadeMux
    port map (
            O => \N__32403\,
            I => \N__32365\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32359\
        );

    \I__7724\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32356\
        );

    \I__7723\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32353\
        );

    \I__7722\ : InMux
    port map (
            O => \N__32395\,
            I => \N__32346\
        );

    \I__7721\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32343\
        );

    \I__7720\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32340\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__32386\,
            I => \N__32335\
        );

    \I__7718\ : IoSpan4Mux
    port map (
            O => \N__32381\,
            I => \N__32335\
        );

    \I__7717\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32332\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__32377\,
            I => \N__32325\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32325\
        );

    \I__7714\ : Span4Mux_s2_h
    port map (
            O => \N__32371\,
            I => \N__32325\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32320\
        );

    \I__7712\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32317\
        );

    \I__7711\ : CascadeMux
    port map (
            O => \N__32364\,
            I => \N__32313\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__32363\,
            I => \N__32310\
        );

    \I__7709\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32307\
        );

    \I__7708\ : Span4Mux_s3_h
    port map (
            O => \N__32359\,
            I => \N__32300\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__32356\,
            I => \N__32300\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__32353\,
            I => \N__32300\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__32352\,
            I => \N__32296\
        );

    \I__7704\ : CascadeMux
    port map (
            O => \N__32351\,
            I => \N__32293\
        );

    \I__7703\ : CascadeMux
    port map (
            O => \N__32350\,
            I => \N__32290\
        );

    \I__7702\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32286\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__32346\,
            I => \N__32279\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32279\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__32340\,
            I => \N__32279\
        );

    \I__7698\ : Span4Mux_s2_h
    port map (
            O => \N__32335\,
            I => \N__32276\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__32332\,
            I => \N__32271\
        );

    \I__7696\ : Span4Mux_h
    port map (
            O => \N__32325\,
            I => \N__32271\
        );

    \I__7695\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32268\
        );

    \I__7694\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32265\
        );

    \I__7693\ : Span4Mux_v
    port map (
            O => \N__32320\,
            I => \N__32259\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__32317\,
            I => \N__32259\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__32316\,
            I => \N__32256\
        );

    \I__7690\ : InMux
    port map (
            O => \N__32313\,
            I => \N__32253\
        );

    \I__7689\ : InMux
    port map (
            O => \N__32310\,
            I => \N__32250\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__32307\,
            I => \N__32245\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__32300\,
            I => \N__32245\
        );

    \I__7686\ : CascadeMux
    port map (
            O => \N__32299\,
            I => \N__32241\
        );

    \I__7685\ : InMux
    port map (
            O => \N__32296\,
            I => \N__32237\
        );

    \I__7684\ : InMux
    port map (
            O => \N__32293\,
            I => \N__32234\
        );

    \I__7683\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32231\
        );

    \I__7682\ : CascadeMux
    port map (
            O => \N__32289\,
            I => \N__32227\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__32286\,
            I => \N__32224\
        );

    \I__7680\ : Span4Mux_v
    port map (
            O => \N__32279\,
            I => \N__32215\
        );

    \I__7679\ : Span4Mux_h
    port map (
            O => \N__32276\,
            I => \N__32215\
        );

    \I__7678\ : Span4Mux_v
    port map (
            O => \N__32271\,
            I => \N__32215\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__32268\,
            I => \N__32215\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32212\
        );

    \I__7675\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32209\
        );

    \I__7674\ : Span4Mux_s2_v
    port map (
            O => \N__32259\,
            I => \N__32206\
        );

    \I__7673\ : InMux
    port map (
            O => \N__32256\,
            I => \N__32203\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__32253\,
            I => \N__32200\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__32250\,
            I => \N__32195\
        );

    \I__7670\ : Span4Mux_v
    port map (
            O => \N__32245\,
            I => \N__32195\
        );

    \I__7669\ : InMux
    port map (
            O => \N__32244\,
            I => \N__32192\
        );

    \I__7668\ : InMux
    port map (
            O => \N__32241\,
            I => \N__32189\
        );

    \I__7667\ : InMux
    port map (
            O => \N__32240\,
            I => \N__32186\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__32237\,
            I => \N__32179\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__32234\,
            I => \N__32179\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__32231\,
            I => \N__32179\
        );

    \I__7663\ : CascadeMux
    port map (
            O => \N__32230\,
            I => \N__32176\
        );

    \I__7662\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32173\
        );

    \I__7661\ : Span4Mux_h
    port map (
            O => \N__32224\,
            I => \N__32168\
        );

    \I__7660\ : Span4Mux_h
    port map (
            O => \N__32215\,
            I => \N__32168\
        );

    \I__7659\ : Span4Mux_h
    port map (
            O => \N__32212\,
            I => \N__32165\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__32209\,
            I => \N__32160\
        );

    \I__7657\ : Span4Mux_h
    port map (
            O => \N__32206\,
            I => \N__32160\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__32203\,
            I => \N__32153\
        );

    \I__7655\ : Span4Mux_s2_v
    port map (
            O => \N__32200\,
            I => \N__32153\
        );

    \I__7654\ : Span4Mux_s3_h
    port map (
            O => \N__32195\,
            I => \N__32153\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__32192\,
            I => \N__32144\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__32189\,
            I => \N__32144\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__32186\,
            I => \N__32144\
        );

    \I__7650\ : Span12Mux_s7_h
    port map (
            O => \N__32179\,
            I => \N__32144\
        );

    \I__7649\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32141\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__32173\,
            I => \N__32136\
        );

    \I__7647\ : Span4Mux_v
    port map (
            O => \N__32168\,
            I => \N__32136\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__32165\,
            I => \processor_zipi8.arith_logical_result_0\
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__32160\,
            I => \processor_zipi8.arith_logical_result_0\
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__32153\,
            I => \processor_zipi8.arith_logical_result_0\
        );

    \I__7643\ : Odrv12
    port map (
            O => \N__32144\,
            I => \processor_zipi8.arith_logical_result_0\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__32141\,
            I => \processor_zipi8.arith_logical_result_0\
        );

    \I__7641\ : Odrv4
    port map (
            O => \N__32136\,
            I => \processor_zipi8.arith_logical_result_0\
        );

    \I__7640\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32116\
        );

    \I__7639\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32112\
        );

    \I__7638\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32106\
        );

    \I__7637\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32103\
        );

    \I__7636\ : CascadeMux
    port map (
            O => \N__32119\,
            I => \N__32094\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__32116\,
            I => \N__32089\
        );

    \I__7634\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32084\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__32112\,
            I => \N__32081\
        );

    \I__7632\ : CascadeMux
    port map (
            O => \N__32111\,
            I => \N__32076\
        );

    \I__7631\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32073\
        );

    \I__7630\ : CascadeMux
    port map (
            O => \N__32109\,
            I => \N__32070\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__32065\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32065\
        );

    \I__7627\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32062\
        );

    \I__7626\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32059\
        );

    \I__7625\ : CascadeMux
    port map (
            O => \N__32100\,
            I => \N__32055\
        );

    \I__7624\ : CascadeMux
    port map (
            O => \N__32099\,
            I => \N__32052\
        );

    \I__7623\ : CascadeMux
    port map (
            O => \N__32098\,
            I => \N__32049\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__32097\,
            I => \N__32046\
        );

    \I__7621\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32043\
        );

    \I__7620\ : InMux
    port map (
            O => \N__32093\,
            I => \N__32040\
        );

    \I__7619\ : InMux
    port map (
            O => \N__32092\,
            I => \N__32037\
        );

    \I__7618\ : Span4Mux_v
    port map (
            O => \N__32089\,
            I => \N__32034\
        );

    \I__7617\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32031\
        );

    \I__7616\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32028\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__32084\,
            I => \N__32019\
        );

    \I__7614\ : Span4Mux_s1_h
    port map (
            O => \N__32081\,
            I => \N__32016\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__32080\,
            I => \N__32013\
        );

    \I__7612\ : InMux
    port map (
            O => \N__32079\,
            I => \N__32010\
        );

    \I__7611\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32007\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__32073\,
            I => \N__32004\
        );

    \I__7609\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32001\
        );

    \I__7608\ : Span4Mux_s3_h
    port map (
            O => \N__32065\,
            I => \N__31998\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__32062\,
            I => \N__31992\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__32059\,
            I => \N__31992\
        );

    \I__7605\ : InMux
    port map (
            O => \N__32058\,
            I => \N__31989\
        );

    \I__7604\ : InMux
    port map (
            O => \N__32055\,
            I => \N__31985\
        );

    \I__7603\ : InMux
    port map (
            O => \N__32052\,
            I => \N__31982\
        );

    \I__7602\ : InMux
    port map (
            O => \N__32049\,
            I => \N__31979\
        );

    \I__7601\ : InMux
    port map (
            O => \N__32046\,
            I => \N__31976\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__31973\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__31968\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__31968\
        );

    \I__7597\ : IoSpan4Mux
    port map (
            O => \N__32034\,
            I => \N__31963\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__32031\,
            I => \N__31963\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__32028\,
            I => \N__31960\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__32027\,
            I => \N__31955\
        );

    \I__7593\ : InMux
    port map (
            O => \N__32026\,
            I => \N__31952\
        );

    \I__7592\ : InMux
    port map (
            O => \N__32025\,
            I => \N__31949\
        );

    \I__7591\ : InMux
    port map (
            O => \N__32024\,
            I => \N__31946\
        );

    \I__7590\ : InMux
    port map (
            O => \N__32023\,
            I => \N__31943\
        );

    \I__7589\ : InMux
    port map (
            O => \N__32022\,
            I => \N__31940\
        );

    \I__7588\ : Span4Mux_s1_h
    port map (
            O => \N__32019\,
            I => \N__31937\
        );

    \I__7587\ : Span4Mux_v
    port map (
            O => \N__32016\,
            I => \N__31934\
        );

    \I__7586\ : InMux
    port map (
            O => \N__32013\,
            I => \N__31931\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__32010\,
            I => \N__31920\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__32007\,
            I => \N__31920\
        );

    \I__7583\ : Span4Mux_s3_h
    port map (
            O => \N__32004\,
            I => \N__31920\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31920\
        );

    \I__7581\ : Span4Mux_v
    port map (
            O => \N__31998\,
            I => \N__31920\
        );

    \I__7580\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31917\
        );

    \I__7579\ : Span4Mux_s3_h
    port map (
            O => \N__31992\,
            I => \N__31914\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31911\
        );

    \I__7577\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31908\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__31985\,
            I => \N__31905\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31898\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31898\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31898\
        );

    \I__7572\ : Span4Mux_v
    port map (
            O => \N__31973\,
            I => \N__31889\
        );

    \I__7571\ : Span4Mux_v
    port map (
            O => \N__31968\,
            I => \N__31889\
        );

    \I__7570\ : Span4Mux_s3_h
    port map (
            O => \N__31963\,
            I => \N__31889\
        );

    \I__7569\ : Span4Mux_s3_h
    port map (
            O => \N__31960\,
            I => \N__31889\
        );

    \I__7568\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31886\
        );

    \I__7567\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31883\
        );

    \I__7566\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31880\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31871\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__31949\,
            I => \N__31871\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__31946\,
            I => \N__31871\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__31943\,
            I => \N__31871\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31868\
        );

    \I__7560\ : Span4Mux_v
    port map (
            O => \N__31937\,
            I => \N__31863\
        );

    \I__7559\ : Span4Mux_v
    port map (
            O => \N__31934\,
            I => \N__31863\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31858\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__31920\,
            I => \N__31858\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__31917\,
            I => \N__31851\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__31914\,
            I => \N__31851\
        );

    \I__7554\ : Span4Mux_s3_h
    port map (
            O => \N__31911\,
            I => \N__31851\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31842\
        );

    \I__7552\ : Span4Mux_h
    port map (
            O => \N__31905\,
            I => \N__31842\
        );

    \I__7551\ : Span4Mux_v
    port map (
            O => \N__31898\,
            I => \N__31842\
        );

    \I__7550\ : Span4Mux_h
    port map (
            O => \N__31889\,
            I => \N__31842\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__31886\,
            I => \N__31832\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__31883\,
            I => \N__31832\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31832\
        );

    \I__7546\ : Span12Mux_v
    port map (
            O => \N__31871\,
            I => \N__31832\
        );

    \I__7545\ : Span4Mux_s2_v
    port map (
            O => \N__31868\,
            I => \N__31827\
        );

    \I__7544\ : Span4Mux_h
    port map (
            O => \N__31863\,
            I => \N__31827\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__31858\,
            I => \N__31824\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__31851\,
            I => \N__31819\
        );

    \I__7541\ : Span4Mux_v
    port map (
            O => \N__31842\,
            I => \N__31819\
        );

    \I__7540\ : InMux
    port map (
            O => \N__31841\,
            I => \N__31816\
        );

    \I__7539\ : Odrv12
    port map (
            O => \N__31832\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197\
        );

    \I__7538\ : Odrv4
    port map (
            O => \N__31827\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197\
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__31824\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197\
        );

    \I__7536\ : Odrv4
    port map (
            O => \N__31819\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__31816\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197\
        );

    \I__7534\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31802\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__31802\,
            I => \N__31798\
        );

    \I__7532\ : InMux
    port map (
            O => \N__31801\,
            I => \N__31795\
        );

    \I__7531\ : Span4Mux_h
    port map (
            O => \N__31798\,
            I => \N__31792\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__31795\,
            I => \N__31789\
        );

    \I__7529\ : Span4Mux_s0_h
    port map (
            O => \N__31792\,
            I => \N__31786\
        );

    \I__7528\ : Span4Mux_h
    port map (
            O => \N__31789\,
            I => \N__31783\
        );

    \I__7527\ : Odrv4
    port map (
            O => \N__31786\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0\
        );

    \I__7526\ : Odrv4
    port map (
            O => \N__31783\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0\
        );

    \I__7525\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31772\
        );

    \I__7524\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31772\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__31772\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_7\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__31769\,
            I => \N__31765\
        );

    \I__7521\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31760\
        );

    \I__7520\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31760\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__31760\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_7\
        );

    \I__7518\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31754\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__31754\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_7\
        );

    \I__7516\ : CascadeMux
    port map (
            O => \N__31751\,
            I => \N__31746\
        );

    \I__7515\ : InMux
    port map (
            O => \N__31750\,
            I => \N__31738\
        );

    \I__7514\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31725\
        );

    \I__7513\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31725\
        );

    \I__7512\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31725\
        );

    \I__7511\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31722\
        );

    \I__7510\ : CascadeMux
    port map (
            O => \N__31743\,
            I => \N__31719\
        );

    \I__7509\ : CascadeMux
    port map (
            O => \N__31742\,
            I => \N__31714\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__31741\,
            I => \N__31709\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__31738\,
            I => \N__31685\
        );

    \I__7506\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31664\
        );

    \I__7505\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31664\
        );

    \I__7504\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31664\
        );

    \I__7503\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31664\
        );

    \I__7502\ : CascadeMux
    port map (
            O => \N__31733\,
            I => \N__31660\
        );

    \I__7501\ : CascadeMux
    port map (
            O => \N__31732\,
            I => \N__31657\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31652\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31652\
        );

    \I__7498\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31647\
        );

    \I__7497\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31647\
        );

    \I__7496\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31642\
        );

    \I__7495\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31642\
        );

    \I__7494\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31639\
        );

    \I__7493\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31632\
        );

    \I__7492\ : InMux
    port map (
            O => \N__31709\,
            I => \N__31632\
        );

    \I__7491\ : InMux
    port map (
            O => \N__31708\,
            I => \N__31632\
        );

    \I__7490\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31625\
        );

    \I__7489\ : InMux
    port map (
            O => \N__31706\,
            I => \N__31625\
        );

    \I__7488\ : InMux
    port map (
            O => \N__31705\,
            I => \N__31625\
        );

    \I__7487\ : CascadeMux
    port map (
            O => \N__31704\,
            I => \N__31620\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__31703\,
            I => \N__31617\
        );

    \I__7485\ : InMux
    port map (
            O => \N__31702\,
            I => \N__31609\
        );

    \I__7484\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31606\
        );

    \I__7483\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31601\
        );

    \I__7482\ : InMux
    port map (
            O => \N__31699\,
            I => \N__31601\
        );

    \I__7481\ : InMux
    port map (
            O => \N__31698\,
            I => \N__31598\
        );

    \I__7480\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31595\
        );

    \I__7479\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31592\
        );

    \I__7478\ : CascadeMux
    port map (
            O => \N__31695\,
            I => \N__31586\
        );

    \I__7477\ : InMux
    port map (
            O => \N__31694\,
            I => \N__31578\
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__31693\,
            I => \N__31565\
        );

    \I__7475\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31558\
        );

    \I__7474\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31558\
        );

    \I__7473\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31558\
        );

    \I__7472\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31553\
        );

    \I__7471\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31553\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__31685\,
            I => \N__31549\
        );

    \I__7469\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31542\
        );

    \I__7468\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31542\
        );

    \I__7467\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31542\
        );

    \I__7466\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31525\
        );

    \I__7465\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31525\
        );

    \I__7464\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31525\
        );

    \I__7463\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31525\
        );

    \I__7462\ : InMux
    port map (
            O => \N__31677\,
            I => \N__31525\
        );

    \I__7461\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31518\
        );

    \I__7460\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31518\
        );

    \I__7459\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31518\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__31673\,
            I => \N__31509\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__31664\,
            I => \N__31504\
        );

    \I__7456\ : InMux
    port map (
            O => \N__31663\,
            I => \N__31497\
        );

    \I__7455\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31497\
        );

    \I__7454\ : InMux
    port map (
            O => \N__31657\,
            I => \N__31497\
        );

    \I__7453\ : Span4Mux_v
    port map (
            O => \N__31652\,
            I => \N__31490\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__31647\,
            I => \N__31490\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__31642\,
            I => \N__31490\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__31639\,
            I => \N__31483\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__31632\,
            I => \N__31483\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__31625\,
            I => \N__31483\
        );

    \I__7447\ : InMux
    port map (
            O => \N__31624\,
            I => \N__31472\
        );

    \I__7446\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31472\
        );

    \I__7445\ : InMux
    port map (
            O => \N__31620\,
            I => \N__31472\
        );

    \I__7444\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31472\
        );

    \I__7443\ : InMux
    port map (
            O => \N__31616\,
            I => \N__31472\
        );

    \I__7442\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31463\
        );

    \I__7441\ : InMux
    port map (
            O => \N__31614\,
            I => \N__31463\
        );

    \I__7440\ : InMux
    port map (
            O => \N__31613\,
            I => \N__31463\
        );

    \I__7439\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31463\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__31609\,
            I => \N__31454\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__31606\,
            I => \N__31454\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__31601\,
            I => \N__31454\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__31598\,
            I => \N__31454\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__31595\,
            I => \N__31449\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__31592\,
            I => \N__31449\
        );

    \I__7432\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31440\
        );

    \I__7431\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31440\
        );

    \I__7430\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31440\
        );

    \I__7429\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31440\
        );

    \I__7428\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31429\
        );

    \I__7427\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31429\
        );

    \I__7426\ : InMux
    port map (
            O => \N__31583\,
            I => \N__31429\
        );

    \I__7425\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31429\
        );

    \I__7424\ : InMux
    port map (
            O => \N__31581\,
            I => \N__31429\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__31578\,
            I => \N__31421\
        );

    \I__7422\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31414\
        );

    \I__7421\ : InMux
    port map (
            O => \N__31576\,
            I => \N__31414\
        );

    \I__7420\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31414\
        );

    \I__7419\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31409\
        );

    \I__7418\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31409\
        );

    \I__7417\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31404\
        );

    \I__7416\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31404\
        );

    \I__7415\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31399\
        );

    \I__7414\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31399\
        );

    \I__7413\ : CascadeMux
    port map (
            O => \N__31568\,
            I => \N__31395\
        );

    \I__7412\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31387\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__31558\,
            I => \N__31381\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__31553\,
            I => \N__31378\
        );

    \I__7409\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31375\
        );

    \I__7408\ : Span4Mux_h
    port map (
            O => \N__31549\,
            I => \N__31370\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__31542\,
            I => \N__31370\
        );

    \I__7406\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31359\
        );

    \I__7405\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31359\
        );

    \I__7404\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31359\
        );

    \I__7403\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31359\
        );

    \I__7402\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31359\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__31536\,
            I => \N__31356\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__31525\,
            I => \N__31353\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__31518\,
            I => \N__31350\
        );

    \I__7398\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31343\
        );

    \I__7397\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31343\
        );

    \I__7396\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31343\
        );

    \I__7395\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31327\
        );

    \I__7394\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31327\
        );

    \I__7393\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31327\
        );

    \I__7392\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31327\
        );

    \I__7391\ : CascadeMux
    port map (
            O => \N__31508\,
            I => \N__31322\
        );

    \I__7390\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31317\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__31504\,
            I => \N__31306\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__31497\,
            I => \N__31306\
        );

    \I__7387\ : Span4Mux_h
    port map (
            O => \N__31490\,
            I => \N__31306\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__31483\,
            I => \N__31306\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__31472\,
            I => \N__31306\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__31463\,
            I => \N__31302\
        );

    \I__7383\ : Span4Mux_v
    port map (
            O => \N__31454\,
            I => \N__31297\
        );

    \I__7382\ : Span4Mux_s1_h
    port map (
            O => \N__31449\,
            I => \N__31297\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__31440\,
            I => \N__31292\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31292\
        );

    \I__7379\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31281\
        );

    \I__7378\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31281\
        );

    \I__7377\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31281\
        );

    \I__7376\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31281\
        );

    \I__7375\ : InMux
    port map (
            O => \N__31424\,
            I => \N__31281\
        );

    \I__7374\ : Span4Mux_v
    port map (
            O => \N__31421\,
            I => \N__31274\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__31414\,
            I => \N__31271\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__31409\,
            I => \N__31264\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31264\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__31399\,
            I => \N__31264\
        );

    \I__7369\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31255\
        );

    \I__7368\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31255\
        );

    \I__7367\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31255\
        );

    \I__7366\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31255\
        );

    \I__7365\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31248\
        );

    \I__7364\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31248\
        );

    \I__7363\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31248\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__31387\,
            I => \N__31245\
        );

    \I__7361\ : InMux
    port map (
            O => \N__31386\,
            I => \N__31238\
        );

    \I__7360\ : InMux
    port map (
            O => \N__31385\,
            I => \N__31238\
        );

    \I__7359\ : InMux
    port map (
            O => \N__31384\,
            I => \N__31238\
        );

    \I__7358\ : Span4Mux_s2_h
    port map (
            O => \N__31381\,
            I => \N__31231\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__31378\,
            I => \N__31231\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31231\
        );

    \I__7355\ : Span4Mux_v
    port map (
            O => \N__31370\,
            I => \N__31228\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__31359\,
            I => \N__31225\
        );

    \I__7353\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31222\
        );

    \I__7352\ : Span4Mux_h
    port map (
            O => \N__31353\,
            I => \N__31210\
        );

    \I__7351\ : Span4Mux_h
    port map (
            O => \N__31350\,
            I => \N__31210\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__31343\,
            I => \N__31210\
        );

    \I__7349\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31195\
        );

    \I__7348\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31195\
        );

    \I__7347\ : InMux
    port map (
            O => \N__31340\,
            I => \N__31195\
        );

    \I__7346\ : InMux
    port map (
            O => \N__31339\,
            I => \N__31195\
        );

    \I__7345\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31195\
        );

    \I__7344\ : InMux
    port map (
            O => \N__31337\,
            I => \N__31195\
        );

    \I__7343\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31195\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__31327\,
            I => \N__31192\
        );

    \I__7341\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31181\
        );

    \I__7340\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31181\
        );

    \I__7339\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31181\
        );

    \I__7338\ : InMux
    port map (
            O => \N__31321\,
            I => \N__31181\
        );

    \I__7337\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31181\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__31317\,
            I => \N__31176\
        );

    \I__7335\ : Span4Mux_h
    port map (
            O => \N__31306\,
            I => \N__31176\
        );

    \I__7334\ : CascadeMux
    port map (
            O => \N__31305\,
            I => \N__31169\
        );

    \I__7333\ : Span4Mux_h
    port map (
            O => \N__31302\,
            I => \N__31166\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__31297\,
            I => \N__31159\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__31292\,
            I => \N__31159\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31159\
        );

    \I__7329\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31150\
        );

    \I__7328\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31150\
        );

    \I__7327\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31150\
        );

    \I__7326\ : InMux
    port map (
            O => \N__31277\,
            I => \N__31150\
        );

    \I__7325\ : Span4Mux_h
    port map (
            O => \N__31274\,
            I => \N__31141\
        );

    \I__7324\ : Span4Mux_v
    port map (
            O => \N__31271\,
            I => \N__31141\
        );

    \I__7323\ : Span4Mux_v
    port map (
            O => \N__31264\,
            I => \N__31141\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__31255\,
            I => \N__31141\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__31248\,
            I => \N__31134\
        );

    \I__7320\ : Span4Mux_v
    port map (
            O => \N__31245\,
            I => \N__31134\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__31238\,
            I => \N__31134\
        );

    \I__7318\ : Sp12to4
    port map (
            O => \N__31231\,
            I => \N__31131\
        );

    \I__7317\ : Span4Mux_h
    port map (
            O => \N__31228\,
            I => \N__31128\
        );

    \I__7316\ : Span4Mux_h
    port map (
            O => \N__31225\,
            I => \N__31123\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__31222\,
            I => \N__31123\
        );

    \I__7314\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31112\
        );

    \I__7313\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31112\
        );

    \I__7312\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31112\
        );

    \I__7311\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31112\
        );

    \I__7310\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31112\
        );

    \I__7309\ : Span4Mux_v
    port map (
            O => \N__31210\,
            I => \N__31107\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__31195\,
            I => \N__31107\
        );

    \I__7307\ : Span4Mux_h
    port map (
            O => \N__31192\,
            I => \N__31100\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__31181\,
            I => \N__31100\
        );

    \I__7305\ : Span4Mux_v
    port map (
            O => \N__31176\,
            I => \N__31100\
        );

    \I__7304\ : InMux
    port map (
            O => \N__31175\,
            I => \N__31089\
        );

    \I__7303\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31089\
        );

    \I__7302\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31089\
        );

    \I__7301\ : InMux
    port map (
            O => \N__31172\,
            I => \N__31089\
        );

    \I__7300\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31089\
        );

    \I__7299\ : Span4Mux_v
    port map (
            O => \N__31166\,
            I => \N__31078\
        );

    \I__7298\ : Span4Mux_h
    port map (
            O => \N__31159\,
            I => \N__31078\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__31150\,
            I => \N__31078\
        );

    \I__7296\ : Span4Mux_h
    port map (
            O => \N__31141\,
            I => \N__31078\
        );

    \I__7295\ : Span4Mux_h
    port map (
            O => \N__31134\,
            I => \N__31078\
        );

    \I__7294\ : Odrv12
    port map (
            O => \N__31131\,
            I => instruction_9
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__31128\,
            I => instruction_9
        );

    \I__7292\ : Odrv4
    port map (
            O => \N__31123\,
            I => instruction_9
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__31112\,
            I => instruction_9
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__31107\,
            I => instruction_9
        );

    \I__7289\ : Odrv4
    port map (
            O => \N__31100\,
            I => instruction_9
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__31089\,
            I => instruction_9
        );

    \I__7287\ : Odrv4
    port map (
            O => \N__31078\,
            I => instruction_9
        );

    \I__7286\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31057\
        );

    \I__7285\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31054\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__31057\,
            I => \N__31049\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__31049\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__31049\,
            I => \N__31046\
        );

    \I__7281\ : Odrv4
    port map (
            O => \N__31046\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_7\
        );

    \I__7280\ : CascadeMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__7279\ : InMux
    port map (
            O => \N__31040\,
            I => \N__31036\
        );

    \I__7278\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31033\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__31036\,
            I => \N__31028\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__31033\,
            I => \N__31028\
        );

    \I__7275\ : Span4Mux_v
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__31025\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_7\
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__31022\,
            I => \N__31018\
        );

    \I__7272\ : InMux
    port map (
            O => \N__31021\,
            I => \N__31010\
        );

    \I__7271\ : InMux
    port map (
            O => \N__31018\,
            I => \N__31001\
        );

    \I__7270\ : CascadeMux
    port map (
            O => \N__31017\,
            I => \N__30997\
        );

    \I__7269\ : CascadeMux
    port map (
            O => \N__31016\,
            I => \N__30994\
        );

    \I__7268\ : CascadeMux
    port map (
            O => \N__31015\,
            I => \N__30990\
        );

    \I__7267\ : CascadeMux
    port map (
            O => \N__31014\,
            I => \N__30987\
        );

    \I__7266\ : InMux
    port map (
            O => \N__31013\,
            I => \N__30976\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__30970\
        );

    \I__7264\ : InMux
    port map (
            O => \N__31009\,
            I => \N__30967\
        );

    \I__7263\ : InMux
    port map (
            O => \N__31008\,
            I => \N__30962\
        );

    \I__7262\ : InMux
    port map (
            O => \N__31007\,
            I => \N__30962\
        );

    \I__7261\ : InMux
    port map (
            O => \N__31006\,
            I => \N__30957\
        );

    \I__7260\ : InMux
    port map (
            O => \N__31005\,
            I => \N__30957\
        );

    \I__7259\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30954\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__31001\,
            I => \N__30951\
        );

    \I__7257\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30946\
        );

    \I__7256\ : InMux
    port map (
            O => \N__30997\,
            I => \N__30946\
        );

    \I__7255\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30939\
        );

    \I__7254\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30936\
        );

    \I__7253\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30933\
        );

    \I__7252\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30928\
        );

    \I__7251\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30923\
        );

    \I__7250\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30923\
        );

    \I__7249\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30918\
        );

    \I__7248\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30911\
        );

    \I__7247\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30911\
        );

    \I__7246\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30904\
        );

    \I__7245\ : InMux
    port map (
            O => \N__30980\,
            I => \N__30904\
        );

    \I__7244\ : CascadeMux
    port map (
            O => \N__30979\,
            I => \N__30901\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__30976\,
            I => \N__30895\
        );

    \I__7242\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30892\
        );

    \I__7241\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30887\
        );

    \I__7240\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30887\
        );

    \I__7239\ : Span4Mux_s2_h
    port map (
            O => \N__30970\,
            I => \N__30882\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__30967\,
            I => \N__30882\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__30962\,
            I => \N__30877\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__30957\,
            I => \N__30877\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__30954\,
            I => \N__30870\
        );

    \I__7234\ : Span4Mux_s3_v
    port map (
            O => \N__30951\,
            I => \N__30870\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__30946\,
            I => \N__30870\
        );

    \I__7232\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30865\
        );

    \I__7231\ : InMux
    port map (
            O => \N__30944\,
            I => \N__30865\
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__30943\,
            I => \N__30861\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__30942\,
            I => \N__30856\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__30939\,
            I => \N__30849\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__30936\,
            I => \N__30849\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__30933\,
            I => \N__30849\
        );

    \I__7225\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30838\
        );

    \I__7224\ : InMux
    port map (
            O => \N__30931\,
            I => \N__30838\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__30928\,
            I => \N__30830\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__30923\,
            I => \N__30827\
        );

    \I__7221\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30824\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__30921\,
            I => \N__30819\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__30918\,
            I => \N__30816\
        );

    \I__7218\ : InMux
    port map (
            O => \N__30917\,
            I => \N__30813\
        );

    \I__7217\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30810\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__30911\,
            I => \N__30807\
        );

    \I__7215\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30802\
        );

    \I__7214\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30802\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__30904\,
            I => \N__30799\
        );

    \I__7212\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30794\
        );

    \I__7211\ : InMux
    port map (
            O => \N__30900\,
            I => \N__30787\
        );

    \I__7210\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30787\
        );

    \I__7209\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30787\
        );

    \I__7208\ : Span4Mux_s3_v
    port map (
            O => \N__30895\,
            I => \N__30780\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__30892\,
            I => \N__30780\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__30887\,
            I => \N__30780\
        );

    \I__7205\ : Span4Mux_h
    port map (
            O => \N__30882\,
            I => \N__30771\
        );

    \I__7204\ : Span4Mux_v
    port map (
            O => \N__30877\,
            I => \N__30771\
        );

    \I__7203\ : Span4Mux_v
    port map (
            O => \N__30870\,
            I => \N__30771\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__30865\,
            I => \N__30771\
        );

    \I__7201\ : InMux
    port map (
            O => \N__30864\,
            I => \N__30768\
        );

    \I__7200\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30765\
        );

    \I__7199\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30760\
        );

    \I__7198\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30760\
        );

    \I__7197\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30757\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__30849\,
            I => \N__30754\
        );

    \I__7195\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30749\
        );

    \I__7194\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30749\
        );

    \I__7193\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30744\
        );

    \I__7192\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30744\
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__30844\,
            I => \N__30741\
        );

    \I__7190\ : CascadeMux
    port map (
            O => \N__30843\,
            I => \N__30738\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30735\
        );

    \I__7188\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30730\
        );

    \I__7187\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30730\
        );

    \I__7186\ : InMux
    port map (
            O => \N__30835\,
            I => \N__30723\
        );

    \I__7185\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30723\
        );

    \I__7184\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30723\
        );

    \I__7183\ : Span4Mux_v
    port map (
            O => \N__30830\,
            I => \N__30716\
        );

    \I__7182\ : Span4Mux_v
    port map (
            O => \N__30827\,
            I => \N__30716\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__30824\,
            I => \N__30716\
        );

    \I__7180\ : InMux
    port map (
            O => \N__30823\,
            I => \N__30709\
        );

    \I__7179\ : InMux
    port map (
            O => \N__30822\,
            I => \N__30709\
        );

    \I__7178\ : InMux
    port map (
            O => \N__30819\,
            I => \N__30709\
        );

    \I__7177\ : Span4Mux_v
    port map (
            O => \N__30816\,
            I => \N__30704\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__30813\,
            I => \N__30704\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__30810\,
            I => \N__30699\
        );

    \I__7174\ : Span4Mux_s3_v
    port map (
            O => \N__30807\,
            I => \N__30699\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__30802\,
            I => \N__30694\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__30799\,
            I => \N__30694\
        );

    \I__7171\ : InMux
    port map (
            O => \N__30798\,
            I => \N__30685\
        );

    \I__7170\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30685\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30682\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__30787\,
            I => \N__30675\
        );

    \I__7167\ : Span4Mux_v
    port map (
            O => \N__30780\,
            I => \N__30675\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__30771\,
            I => \N__30675\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__30768\,
            I => \N__30670\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30670\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__30760\,
            I => \N__30667\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__30757\,
            I => \N__30660\
        );

    \I__7161\ : Span4Mux_h
    port map (
            O => \N__30754\,
            I => \N__30660\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__30749\,
            I => \N__30660\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__30744\,
            I => \N__30653\
        );

    \I__7158\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30648\
        );

    \I__7157\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30648\
        );

    \I__7156\ : Span4Mux_v
    port map (
            O => \N__30735\,
            I => \N__30637\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__30730\,
            I => \N__30637\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__30723\,
            I => \N__30637\
        );

    \I__7153\ : Span4Mux_h
    port map (
            O => \N__30716\,
            I => \N__30637\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__30709\,
            I => \N__30637\
        );

    \I__7151\ : Span4Mux_h
    port map (
            O => \N__30704\,
            I => \N__30628\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__30699\,
            I => \N__30628\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__30694\,
            I => \N__30628\
        );

    \I__7148\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30623\
        );

    \I__7147\ : InMux
    port map (
            O => \N__30692\,
            I => \N__30623\
        );

    \I__7146\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30618\
        );

    \I__7145\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30618\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__30685\,
            I => \N__30609\
        );

    \I__7143\ : Span4Mux_v
    port map (
            O => \N__30682\,
            I => \N__30609\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__30675\,
            I => \N__30609\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__30670\,
            I => \N__30609\
        );

    \I__7140\ : Span4Mux_s2_h
    port map (
            O => \N__30667\,
            I => \N__30604\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__30660\,
            I => \N__30604\
        );

    \I__7138\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30595\
        );

    \I__7137\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30595\
        );

    \I__7136\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30595\
        );

    \I__7135\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30595\
        );

    \I__7134\ : Span4Mux_v
    port map (
            O => \N__30653\,
            I => \N__30588\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__30648\,
            I => \N__30588\
        );

    \I__7132\ : Span4Mux_h
    port map (
            O => \N__30637\,
            I => \N__30588\
        );

    \I__7131\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30583\
        );

    \I__7130\ : InMux
    port map (
            O => \N__30635\,
            I => \N__30583\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__30628\,
            I => instruction_8
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__30623\,
            I => instruction_8
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__30618\,
            I => instruction_8
        );

    \I__7126\ : Odrv4
    port map (
            O => \N__30609\,
            I => instruction_8
        );

    \I__7125\ : Odrv4
    port map (
            O => \N__30604\,
            I => instruction_8
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__30595\,
            I => instruction_8
        );

    \I__7123\ : Odrv4
    port map (
            O => \N__30588\,
            I => instruction_8
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__30583\,
            I => instruction_8
        );

    \I__7121\ : InMux
    port map (
            O => \N__30566\,
            I => \N__30563\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__30563\,
            I => \N__30560\
        );

    \I__7119\ : Odrv12
    port map (
            O => \N__30560\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_7\
        );

    \I__7118\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30554\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__30554\,
            I => \N__30550\
        );

    \I__7116\ : InMux
    port map (
            O => \N__30553\,
            I => \N__30547\
        );

    \I__7115\ : Span4Mux_v
    port map (
            O => \N__30550\,
            I => \N__30544\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__30547\,
            I => \N__30541\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__30544\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0\
        );

    \I__7112\ : Odrv12
    port map (
            O => \N__30541\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0\
        );

    \I__7111\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30532\
        );

    \I__7110\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30529\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__30532\,
            I => \N__30524\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30524\
        );

    \I__7107\ : Span4Mux_v
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__30521\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_3\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__30518\,
            I => \N__30515\
        );

    \I__7104\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30511\
        );

    \I__7103\ : CascadeMux
    port map (
            O => \N__30514\,
            I => \N__30504\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__30511\,
            I => \N__30501\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__30510\,
            I => \N__30495\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__30509\,
            I => \N__30486\
        );

    \I__7099\ : CascadeMux
    port map (
            O => \N__30508\,
            I => \N__30482\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__30507\,
            I => \N__30478\
        );

    \I__7097\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30474\
        );

    \I__7096\ : Span4Mux_s2_h
    port map (
            O => \N__30501\,
            I => \N__30468\
        );

    \I__7095\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30465\
        );

    \I__7094\ : CascadeMux
    port map (
            O => \N__30499\,
            I => \N__30458\
        );

    \I__7093\ : CascadeMux
    port map (
            O => \N__30498\,
            I => \N__30455\
        );

    \I__7092\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30452\
        );

    \I__7091\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30449\
        );

    \I__7090\ : InMux
    port map (
            O => \N__30493\,
            I => \N__30445\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__30492\,
            I => \N__30441\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__30491\,
            I => \N__30436\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__30490\,
            I => \N__30433\
        );

    \I__7086\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30430\
        );

    \I__7085\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30427\
        );

    \I__7084\ : InMux
    port map (
            O => \N__30485\,
            I => \N__30424\
        );

    \I__7083\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30421\
        );

    \I__7082\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30418\
        );

    \I__7081\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30415\
        );

    \I__7080\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30412\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30409\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__30473\,
            I => \N__30406\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__30472\,
            I => \N__30403\
        );

    \I__7076\ : CascadeMux
    port map (
            O => \N__30471\,
            I => \N__30400\
        );

    \I__7075\ : Span4Mux_v
    port map (
            O => \N__30468\,
            I => \N__30395\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__30465\,
            I => \N__30395\
        );

    \I__7073\ : InMux
    port map (
            O => \N__30464\,
            I => \N__30391\
        );

    \I__7072\ : CascadeMux
    port map (
            O => \N__30463\,
            I => \N__30387\
        );

    \I__7071\ : CascadeMux
    port map (
            O => \N__30462\,
            I => \N__30383\
        );

    \I__7070\ : InMux
    port map (
            O => \N__30461\,
            I => \N__30380\
        );

    \I__7069\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30377\
        );

    \I__7068\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30374\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__30452\,
            I => \N__30371\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__30449\,
            I => \N__30368\
        );

    \I__7065\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30365\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__30445\,
            I => \N__30362\
        );

    \I__7063\ : CascadeMux
    port map (
            O => \N__30444\,
            I => \N__30359\
        );

    \I__7062\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30356\
        );

    \I__7061\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30353\
        );

    \I__7060\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30350\
        );

    \I__7059\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30347\
        );

    \I__7058\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30344\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__30430\,
            I => \N__30341\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__30427\,
            I => \N__30338\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30335\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__30421\,
            I => \N__30332\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30323\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__30415\,
            I => \N__30323\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__30412\,
            I => \N__30323\
        );

    \I__7050\ : Span4Mux_v
    port map (
            O => \N__30409\,
            I => \N__30323\
        );

    \I__7049\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30320\
        );

    \I__7048\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30317\
        );

    \I__7047\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30314\
        );

    \I__7046\ : Span4Mux_h
    port map (
            O => \N__30395\,
            I => \N__30311\
        );

    \I__7045\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30308\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__30391\,
            I => \N__30305\
        );

    \I__7043\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30302\
        );

    \I__7042\ : InMux
    port map (
            O => \N__30387\,
            I => \N__30299\
        );

    \I__7041\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30296\
        );

    \I__7040\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30293\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__30380\,
            I => \N__30288\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__30377\,
            I => \N__30288\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__30374\,
            I => \N__30281\
        );

    \I__7036\ : Span4Mux_v
    port map (
            O => \N__30371\,
            I => \N__30281\
        );

    \I__7035\ : Span4Mux_v
    port map (
            O => \N__30368\,
            I => \N__30281\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__30365\,
            I => \N__30276\
        );

    \I__7033\ : Span4Mux_s3_v
    port map (
            O => \N__30362\,
            I => \N__30276\
        );

    \I__7032\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30273\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__30356\,
            I => \N__30270\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30254\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__30350\,
            I => \N__30254\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30254\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__30344\,
            I => \N__30254\
        );

    \I__7026\ : Span4Mux_v
    port map (
            O => \N__30341\,
            I => \N__30254\
        );

    \I__7025\ : Span4Mux_h
    port map (
            O => \N__30338\,
            I => \N__30254\
        );

    \I__7024\ : Span4Mux_s2_v
    port map (
            O => \N__30335\,
            I => \N__30254\
        );

    \I__7023\ : Span4Mux_s3_h
    port map (
            O => \N__30332\,
            I => \N__30251\
        );

    \I__7022\ : Span4Mux_v
    port map (
            O => \N__30323\,
            I => \N__30248\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__30320\,
            I => \N__30241\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__30317\,
            I => \N__30241\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__30314\,
            I => \N__30241\
        );

    \I__7018\ : Sp12to4
    port map (
            O => \N__30311\,
            I => \N__30238\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__30308\,
            I => \N__30235\
        );

    \I__7016\ : Span4Mux_s2_v
    port map (
            O => \N__30305\,
            I => \N__30232\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__30302\,
            I => \N__30229\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__30299\,
            I => \N__30224\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__30296\,
            I => \N__30224\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30219\
        );

    \I__7011\ : Span4Mux_v
    port map (
            O => \N__30288\,
            I => \N__30219\
        );

    \I__7010\ : Span4Mux_v
    port map (
            O => \N__30281\,
            I => \N__30214\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__30276\,
            I => \N__30214\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__30273\,
            I => \N__30211\
        );

    \I__7007\ : Span4Mux_s2_h
    port map (
            O => \N__30270\,
            I => \N__30208\
        );

    \I__7006\ : InMux
    port map (
            O => \N__30269\,
            I => \N__30204\
        );

    \I__7005\ : Span4Mux_v
    port map (
            O => \N__30254\,
            I => \N__30197\
        );

    \I__7004\ : Span4Mux_v
    port map (
            O => \N__30251\,
            I => \N__30197\
        );

    \I__7003\ : Span4Mux_h
    port map (
            O => \N__30248\,
            I => \N__30197\
        );

    \I__7002\ : Span12Mux_s6_h
    port map (
            O => \N__30241\,
            I => \N__30192\
        );

    \I__7001\ : Span12Mux_s3_v
    port map (
            O => \N__30238\,
            I => \N__30192\
        );

    \I__7000\ : Span4Mux_h
    port map (
            O => \N__30235\,
            I => \N__30187\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__30232\,
            I => \N__30187\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__30229\,
            I => \N__30178\
        );

    \I__6997\ : Span4Mux_v
    port map (
            O => \N__30224\,
            I => \N__30178\
        );

    \I__6996\ : Span4Mux_h
    port map (
            O => \N__30219\,
            I => \N__30178\
        );

    \I__6995\ : Span4Mux_h
    port map (
            O => \N__30214\,
            I => \N__30178\
        );

    \I__6994\ : Span4Mux_v
    port map (
            O => \N__30211\,
            I => \N__30173\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__30208\,
            I => \N__30173\
        );

    \I__6992\ : InMux
    port map (
            O => \N__30207\,
            I => \N__30170\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__30204\,
            I => \processor_zipi8.arith_logical_result_5\
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__30197\,
            I => \processor_zipi8.arith_logical_result_5\
        );

    \I__6989\ : Odrv12
    port map (
            O => \N__30192\,
            I => \processor_zipi8.arith_logical_result_5\
        );

    \I__6988\ : Odrv4
    port map (
            O => \N__30187\,
            I => \processor_zipi8.arith_logical_result_5\
        );

    \I__6987\ : Odrv4
    port map (
            O => \N__30178\,
            I => \processor_zipi8.arith_logical_result_5\
        );

    \I__6986\ : Odrv4
    port map (
            O => \N__30173\,
            I => \processor_zipi8.arith_logical_result_5\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__30170\,
            I => \processor_zipi8.arith_logical_result_5\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__30155\,
            I => \N__30151\
        );

    \I__6983\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30141\
        );

    \I__6982\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30138\
        );

    \I__6981\ : CascadeMux
    port map (
            O => \N__30150\,
            I => \N__30131\
        );

    \I__6980\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30128\
        );

    \I__6979\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30125\
        );

    \I__6978\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30122\
        );

    \I__6977\ : CascadeMux
    port map (
            O => \N__30146\,
            I => \N__30118\
        );

    \I__6976\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30112\
        );

    \I__6975\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30109\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__30141\,
            I => \N__30106\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__30138\,
            I => \N__30103\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__30137\,
            I => \N__30100\
        );

    \I__6971\ : CascadeMux
    port map (
            O => \N__30136\,
            I => \N__30097\
        );

    \I__6970\ : CascadeMux
    port map (
            O => \N__30135\,
            I => \N__30094\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__30134\,
            I => \N__30091\
        );

    \I__6968\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30085\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__30128\,
            I => \N__30082\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__30125\,
            I => \N__30077\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__30122\,
            I => \N__30077\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__30121\,
            I => \N__30073\
        );

    \I__6963\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30070\
        );

    \I__6962\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30064\
        );

    \I__6961\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30061\
        );

    \I__6960\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30058\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30048\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__30109\,
            I => \N__30048\
        );

    \I__6957\ : Span4Mux_s2_h
    port map (
            O => \N__30106\,
            I => \N__30048\
        );

    \I__6956\ : Span4Mux_s3_v
    port map (
            O => \N__30103\,
            I => \N__30048\
        );

    \I__6955\ : InMux
    port map (
            O => \N__30100\,
            I => \N__30045\
        );

    \I__6954\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30041\
        );

    \I__6953\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30038\
        );

    \I__6952\ : InMux
    port map (
            O => \N__30091\,
            I => \N__30035\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__30090\,
            I => \N__30031\
        );

    \I__6950\ : InMux
    port map (
            O => \N__30089\,
            I => \N__30028\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__30088\,
            I => \N__30025\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__30085\,
            I => \N__30021\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__30082\,
            I => \N__30016\
        );

    \I__6946\ : Span4Mux_v
    port map (
            O => \N__30077\,
            I => \N__30016\
        );

    \I__6945\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30013\
        );

    \I__6944\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30010\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__30070\,
            I => \N__30007\
        );

    \I__6942\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30004\
        );

    \I__6941\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30001\
        );

    \I__6940\ : InMux
    port map (
            O => \N__30067\,
            I => \N__29998\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__30064\,
            I => \N__29993\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__30061\,
            I => \N__29993\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__30058\,
            I => \N__29990\
        );

    \I__6936\ : InMux
    port map (
            O => \N__30057\,
            I => \N__29987\
        );

    \I__6935\ : Span4Mux_h
    port map (
            O => \N__30048\,
            I => \N__29982\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__30045\,
            I => \N__29982\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__30044\,
            I => \N__29979\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__30041\,
            I => \N__29974\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__30038\,
            I => \N__29974\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__30035\,
            I => \N__29971\
        );

    \I__6929\ : InMux
    port map (
            O => \N__30034\,
            I => \N__29968\
        );

    \I__6928\ : InMux
    port map (
            O => \N__30031\,
            I => \N__29965\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__30028\,
            I => \N__29962\
        );

    \I__6926\ : InMux
    port map (
            O => \N__30025\,
            I => \N__29959\
        );

    \I__6925\ : InMux
    port map (
            O => \N__30024\,
            I => \N__29956\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__30021\,
            I => \N__29953\
        );

    \I__6923\ : Span4Mux_s0_h
    port map (
            O => \N__30016\,
            I => \N__29947\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__30013\,
            I => \N__29944\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__30010\,
            I => \N__29937\
        );

    \I__6920\ : Span4Mux_s3_v
    port map (
            O => \N__30007\,
            I => \N__29937\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__30004\,
            I => \N__29937\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__30001\,
            I => \N__29928\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__29998\,
            I => \N__29928\
        );

    \I__6916\ : Span4Mux_v
    port map (
            O => \N__29993\,
            I => \N__29928\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__29990\,
            I => \N__29928\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__29987\,
            I => \N__29923\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__29982\,
            I => \N__29923\
        );

    \I__6912\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29920\
        );

    \I__6911\ : Span4Mux_s1_h
    port map (
            O => \N__29974\,
            I => \N__29917\
        );

    \I__6910\ : Span4Mux_s2_v
    port map (
            O => \N__29971\,
            I => \N__29914\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__29968\,
            I => \N__29911\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__29965\,
            I => \N__29908\
        );

    \I__6907\ : Span4Mux_h
    port map (
            O => \N__29962\,
            I => \N__29901\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__29959\,
            I => \N__29901\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__29956\,
            I => \N__29901\
        );

    \I__6904\ : Span4Mux_h
    port map (
            O => \N__29953\,
            I => \N__29898\
        );

    \I__6903\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29895\
        );

    \I__6902\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29891\
        );

    \I__6901\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29888\
        );

    \I__6900\ : Span4Mux_h
    port map (
            O => \N__29947\,
            I => \N__29885\
        );

    \I__6899\ : Span4Mux_v
    port map (
            O => \N__29944\,
            I => \N__29878\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__29937\,
            I => \N__29878\
        );

    \I__6897\ : Span4Mux_v
    port map (
            O => \N__29928\,
            I => \N__29878\
        );

    \I__6896\ : Span4Mux_h
    port map (
            O => \N__29923\,
            I => \N__29875\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__29920\,
            I => \N__29866\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__29917\,
            I => \N__29866\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__29914\,
            I => \N__29866\
        );

    \I__6892\ : Span4Mux_v
    port map (
            O => \N__29911\,
            I => \N__29866\
        );

    \I__6891\ : Span4Mux_h
    port map (
            O => \N__29908\,
            I => \N__29861\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__29901\,
            I => \N__29861\
        );

    \I__6889\ : Span4Mux_h
    port map (
            O => \N__29898\,
            I => \N__29856\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__29895\,
            I => \N__29856\
        );

    \I__6887\ : InMux
    port map (
            O => \N__29894\,
            I => \N__29853\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__29891\,
            I => \N__29848\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29848\
        );

    \I__6884\ : Span4Mux_h
    port map (
            O => \N__29885\,
            I => \N__29845\
        );

    \I__6883\ : Sp12to4
    port map (
            O => \N__29878\,
            I => \N__29842\
        );

    \I__6882\ : Span4Mux_s1_h
    port map (
            O => \N__29875\,
            I => \N__29839\
        );

    \I__6881\ : Span4Mux_h
    port map (
            O => \N__29866\,
            I => \N__29834\
        );

    \I__6880\ : Span4Mux_h
    port map (
            O => \N__29861\,
            I => \N__29834\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__29856\,
            I => \N__29831\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__29853\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__29848\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__29845\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\
        );

    \I__6875\ : Odrv12
    port map (
            O => \N__29842\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__29839\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\
        );

    \I__6873\ : Odrv4
    port map (
            O => \N__29834\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\
        );

    \I__6872\ : Odrv4
    port map (
            O => \N__29831\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__29816\,
            I => \N__29813\
        );

    \I__6870\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29809\
        );

    \I__6869\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29806\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__29809\,
            I => \N__29803\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29800\
        );

    \I__6866\ : Span4Mux_v
    port map (
            O => \N__29803\,
            I => \N__29797\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__29800\,
            I => \N__29794\
        );

    \I__6864\ : Span4Mux_h
    port map (
            O => \N__29797\,
            I => \N__29791\
        );

    \I__6863\ : Sp12to4
    port map (
            O => \N__29794\,
            I => \N__29788\
        );

    \I__6862\ : Odrv4
    port map (
            O => \N__29791\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5\
        );

    \I__6861\ : Odrv12
    port map (
            O => \N__29788\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__29783\,
            I => \N__29777\
        );

    \I__6859\ : CascadeMux
    port map (
            O => \N__29782\,
            I => \N__29774\
        );

    \I__6858\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29765\
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__29780\,
            I => \N__29761\
        );

    \I__6856\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29758\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29755\
        );

    \I__6854\ : CascadeMux
    port map (
            O => \N__29773\,
            I => \N__29752\
        );

    \I__6853\ : InMux
    port map (
            O => \N__29772\,
            I => \N__29748\
        );

    \I__6852\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29745\
        );

    \I__6851\ : CascadeMux
    port map (
            O => \N__29770\,
            I => \N__29740\
        );

    \I__6850\ : CascadeMux
    port map (
            O => \N__29769\,
            I => \N__29737\
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__29768\,
            I => \N__29732\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__29765\,
            I => \N__29729\
        );

    \I__6847\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29726\
        );

    \I__6846\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29723\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__29758\,
            I => \N__29717\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29717\
        );

    \I__6843\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29714\
        );

    \I__6842\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29711\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__29748\,
            I => \N__29701\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__29745\,
            I => \N__29698\
        );

    \I__6839\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29695\
        );

    \I__6838\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29692\
        );

    \I__6837\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29688\
        );

    \I__6836\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29685\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__29736\,
            I => \N__29681\
        );

    \I__6834\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29678\
        );

    \I__6833\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29672\
        );

    \I__6832\ : Span4Mux_s3_v
    port map (
            O => \N__29729\,
            I => \N__29665\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29665\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29665\
        );

    \I__6829\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29662\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__29717\,
            I => \N__29659\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__29714\,
            I => \N__29656\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29653\
        );

    \I__6825\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29650\
        );

    \I__6824\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29647\
        );

    \I__6823\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29644\
        );

    \I__6822\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29639\
        );

    \I__6821\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29636\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__29705\,
            I => \N__29633\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__29704\,
            I => \N__29630\
        );

    \I__6818\ : Span4Mux_s2_h
    port map (
            O => \N__29701\,
            I => \N__29621\
        );

    \I__6817\ : Span4Mux_s3_v
    port map (
            O => \N__29698\,
            I => \N__29621\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29621\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__29692\,
            I => \N__29621\
        );

    \I__6814\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29618\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__29688\,
            I => \N__29615\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__29685\,
            I => \N__29612\
        );

    \I__6811\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29609\
        );

    \I__6810\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29606\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__29678\,
            I => \N__29603\
        );

    \I__6808\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29600\
        );

    \I__6807\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29597\
        );

    \I__6806\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29594\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__29672\,
            I => \N__29591\
        );

    \I__6804\ : Span4Mux_v
    port map (
            O => \N__29665\,
            I => \N__29586\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__29662\,
            I => \N__29586\
        );

    \I__6802\ : Span4Mux_v
    port map (
            O => \N__29659\,
            I => \N__29581\
        );

    \I__6801\ : Span4Mux_s3_v
    port map (
            O => \N__29656\,
            I => \N__29581\
        );

    \I__6800\ : Span4Mux_s0_h
    port map (
            O => \N__29653\,
            I => \N__29572\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__29650\,
            I => \N__29572\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__29647\,
            I => \N__29572\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__29644\,
            I => \N__29572\
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__29643\,
            I => \N__29569\
        );

    \I__6795\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29566\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__29639\,
            I => \N__29561\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__29636\,
            I => \N__29561\
        );

    \I__6792\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29558\
        );

    \I__6791\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29555\
        );

    \I__6790\ : Span4Mux_h
    port map (
            O => \N__29621\,
            I => \N__29548\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__29618\,
            I => \N__29548\
        );

    \I__6788\ : Span4Mux_v
    port map (
            O => \N__29615\,
            I => \N__29541\
        );

    \I__6787\ : Span4Mux_v
    port map (
            O => \N__29612\,
            I => \N__29541\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__29609\,
            I => \N__29541\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__29606\,
            I => \N__29538\
        );

    \I__6784\ : Span4Mux_h
    port map (
            O => \N__29603\,
            I => \N__29529\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__29600\,
            I => \N__29529\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__29597\,
            I => \N__29529\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__29594\,
            I => \N__29529\
        );

    \I__6780\ : Span4Mux_s3_h
    port map (
            O => \N__29591\,
            I => \N__29524\
        );

    \I__6779\ : Span4Mux_v
    port map (
            O => \N__29586\,
            I => \N__29524\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__29581\,
            I => \N__29519\
        );

    \I__6777\ : Span4Mux_v
    port map (
            O => \N__29572\,
            I => \N__29519\
        );

    \I__6776\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29516\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__29566\,
            I => \N__29513\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__29561\,
            I => \N__29506\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__29558\,
            I => \N__29506\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__29555\,
            I => \N__29506\
        );

    \I__6771\ : InMux
    port map (
            O => \N__29554\,
            I => \N__29503\
        );

    \I__6770\ : InMux
    port map (
            O => \N__29553\,
            I => \N__29500\
        );

    \I__6769\ : Span4Mux_h
    port map (
            O => \N__29548\,
            I => \N__29496\
        );

    \I__6768\ : Span4Mux_h
    port map (
            O => \N__29541\,
            I => \N__29493\
        );

    \I__6767\ : Span4Mux_v
    port map (
            O => \N__29538\,
            I => \N__29490\
        );

    \I__6766\ : Span4Mux_v
    port map (
            O => \N__29529\,
            I => \N__29485\
        );

    \I__6765\ : Span4Mux_h
    port map (
            O => \N__29524\,
            I => \N__29485\
        );

    \I__6764\ : Sp12to4
    port map (
            O => \N__29519\,
            I => \N__29480\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__29516\,
            I => \N__29480\
        );

    \I__6762\ : Span4Mux_h
    port map (
            O => \N__29513\,
            I => \N__29477\
        );

    \I__6761\ : Span4Mux_h
    port map (
            O => \N__29506\,
            I => \N__29470\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29470\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__29500\,
            I => \N__29470\
        );

    \I__6758\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29467\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__29496\,
            I => \N__29460\
        );

    \I__6756\ : Span4Mux_h
    port map (
            O => \N__29493\,
            I => \N__29460\
        );

    \I__6755\ : Span4Mux_h
    port map (
            O => \N__29490\,
            I => \N__29460\
        );

    \I__6754\ : Odrv4
    port map (
            O => \N__29485\,
            I => \processor_zipi8.arith_logical_result_6\
        );

    \I__6753\ : Odrv12
    port map (
            O => \N__29480\,
            I => \processor_zipi8.arith_logical_result_6\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__29477\,
            I => \processor_zipi8.arith_logical_result_6\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__29470\,
            I => \processor_zipi8.arith_logical_result_6\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__29467\,
            I => \processor_zipi8.arith_logical_result_6\
        );

    \I__6749\ : Odrv4
    port map (
            O => \N__29460\,
            I => \processor_zipi8.arith_logical_result_6\
        );

    \I__6748\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29442\
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__29446\,
            I => \N__29439\
        );

    \I__6746\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29434\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29431\
        );

    \I__6744\ : InMux
    port map (
            O => \N__29439\,
            I => \N__29428\
        );

    \I__6743\ : InMux
    port map (
            O => \N__29438\,
            I => \N__29425\
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__29437\,
            I => \N__29422\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__29434\,
            I => \N__29415\
        );

    \I__6740\ : Span4Mux_s1_v
    port map (
            O => \N__29431\,
            I => \N__29415\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__29428\,
            I => \N__29415\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__29425\,
            I => \N__29412\
        );

    \I__6737\ : InMux
    port map (
            O => \N__29422\,
            I => \N__29409\
        );

    \I__6736\ : Span4Mux_h
    port map (
            O => \N__29415\,
            I => \N__29399\
        );

    \I__6735\ : Span4Mux_v
    port map (
            O => \N__29412\,
            I => \N__29399\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29399\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__29408\,
            I => \N__29390\
        );

    \I__6732\ : CascadeMux
    port map (
            O => \N__29407\,
            I => \N__29387\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__29406\,
            I => \N__29384\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__29399\,
            I => \N__29381\
        );

    \I__6729\ : InMux
    port map (
            O => \N__29398\,
            I => \N__29378\
        );

    \I__6728\ : CascadeMux
    port map (
            O => \N__29397\,
            I => \N__29375\
        );

    \I__6727\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29372\
        );

    \I__6726\ : CascadeMux
    port map (
            O => \N__29395\,
            I => \N__29361\
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__29394\,
            I => \N__29358\
        );

    \I__6724\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29353\
        );

    \I__6723\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29350\
        );

    \I__6722\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29347\
        );

    \I__6721\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29344\
        );

    \I__6720\ : Span4Mux_s0_h
    port map (
            O => \N__29381\,
            I => \N__29339\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__29378\,
            I => \N__29339\
        );

    \I__6718\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29336\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__29372\,
            I => \N__29333\
        );

    \I__6716\ : InMux
    port map (
            O => \N__29371\,
            I => \N__29330\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__29370\,
            I => \N__29326\
        );

    \I__6714\ : CascadeMux
    port map (
            O => \N__29369\,
            I => \N__29323\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__29368\,
            I => \N__29320\
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__29367\,
            I => \N__29317\
        );

    \I__6711\ : CascadeMux
    port map (
            O => \N__29366\,
            I => \N__29312\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__29365\,
            I => \N__29308\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__29364\,
            I => \N__29305\
        );

    \I__6708\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29302\
        );

    \I__6707\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29298\
        );

    \I__6706\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29295\
        );

    \I__6705\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29292\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__29353\,
            I => \N__29284\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__29350\,
            I => \N__29284\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__29347\,
            I => \N__29284\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__29344\,
            I => \N__29281\
        );

    \I__6700\ : Span4Mux_v
    port map (
            O => \N__29339\,
            I => \N__29278\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__29336\,
            I => \N__29275\
        );

    \I__6698\ : Span4Mux_s2_v
    port map (
            O => \N__29333\,
            I => \N__29272\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__29330\,
            I => \N__29269\
        );

    \I__6696\ : CascadeMux
    port map (
            O => \N__29329\,
            I => \N__29266\
        );

    \I__6695\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29262\
        );

    \I__6694\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29259\
        );

    \I__6693\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29256\
        );

    \I__6692\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29253\
        );

    \I__6691\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29250\
        );

    \I__6690\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29247\
        );

    \I__6689\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29244\
        );

    \I__6688\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29241\
        );

    \I__6687\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29238\
        );

    \I__6686\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29235\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__29302\,
            I => \N__29232\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__29301\,
            I => \N__29229\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__29298\,
            I => \N__29226\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__29295\,
            I => \N__29223\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__29292\,
            I => \N__29220\
        );

    \I__6680\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29217\
        );

    \I__6679\ : Span4Mux_v
    port map (
            O => \N__29284\,
            I => \N__29214\
        );

    \I__6678\ : Span4Mux_v
    port map (
            O => \N__29281\,
            I => \N__29209\
        );

    \I__6677\ : Span4Mux_h
    port map (
            O => \N__29278\,
            I => \N__29209\
        );

    \I__6676\ : Span4Mux_h
    port map (
            O => \N__29275\,
            I => \N__29202\
        );

    \I__6675\ : Span4Mux_h
    port map (
            O => \N__29272\,
            I => \N__29202\
        );

    \I__6674\ : Span4Mux_s3_h
    port map (
            O => \N__29269\,
            I => \N__29202\
        );

    \I__6673\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29198\
        );

    \I__6672\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29195\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29188\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__29259\,
            I => \N__29188\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29188\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29185\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__29250\,
            I => \N__29176\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__29247\,
            I => \N__29176\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__29244\,
            I => \N__29176\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__29241\,
            I => \N__29176\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__29238\,
            I => \N__29173\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29168\
        );

    \I__6661\ : Span4Mux_h
    port map (
            O => \N__29232\,
            I => \N__29168\
        );

    \I__6660\ : InMux
    port map (
            O => \N__29229\,
            I => \N__29165\
        );

    \I__6659\ : Span4Mux_s3_h
    port map (
            O => \N__29226\,
            I => \N__29158\
        );

    \I__6658\ : Span4Mux_v
    port map (
            O => \N__29223\,
            I => \N__29158\
        );

    \I__6657\ : Span4Mux_v
    port map (
            O => \N__29220\,
            I => \N__29158\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__29217\,
            I => \N__29155\
        );

    \I__6655\ : Span4Mux_h
    port map (
            O => \N__29214\,
            I => \N__29148\
        );

    \I__6654\ : Span4Mux_h
    port map (
            O => \N__29209\,
            I => \N__29148\
        );

    \I__6653\ : Span4Mux_v
    port map (
            O => \N__29202\,
            I => \N__29148\
        );

    \I__6652\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29145\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__29198\,
            I => \N__29142\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29137\
        );

    \I__6649\ : Span12Mux_s5_h
    port map (
            O => \N__29188\,
            I => \N__29137\
        );

    \I__6648\ : Span4Mux_s3_v
    port map (
            O => \N__29185\,
            I => \N__29132\
        );

    \I__6647\ : Span4Mux_v
    port map (
            O => \N__29176\,
            I => \N__29132\
        );

    \I__6646\ : Span4Mux_s3_h
    port map (
            O => \N__29173\,
            I => \N__29127\
        );

    \I__6645\ : Span4Mux_h
    port map (
            O => \N__29168\,
            I => \N__29127\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__29165\,
            I => \N__29122\
        );

    \I__6643\ : Span4Mux_h
    port map (
            O => \N__29158\,
            I => \N__29122\
        );

    \I__6642\ : Span4Mux_h
    port map (
            O => \N__29155\,
            I => \N__29117\
        );

    \I__6641\ : Span4Mux_v
    port map (
            O => \N__29148\,
            I => \N__29117\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__29145\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\
        );

    \I__6639\ : Odrv4
    port map (
            O => \N__29142\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\
        );

    \I__6638\ : Odrv12
    port map (
            O => \N__29137\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__29132\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__29127\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\
        );

    \I__6635\ : Odrv4
    port map (
            O => \N__29122\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\
        );

    \I__6634\ : Odrv4
    port map (
            O => \N__29117\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\
        );

    \I__6633\ : CascadeMux
    port map (
            O => \N__29102\,
            I => \N__29099\
        );

    \I__6632\ : InMux
    port map (
            O => \N__29099\,
            I => \N__29096\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__29096\,
            I => \N__29092\
        );

    \I__6630\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29089\
        );

    \I__6629\ : Span4Mux_s3_v
    port map (
            O => \N__29092\,
            I => \N__29084\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29084\
        );

    \I__6627\ : Span4Mux_v
    port map (
            O => \N__29084\,
            I => \N__29081\
        );

    \I__6626\ : Span4Mux_h
    port map (
            O => \N__29081\,
            I => \N__29078\
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__29078\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_6\
        );

    \I__6624\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29072\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__29072\,
            I => \N__29068\
        );

    \I__6622\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29065\
        );

    \I__6621\ : Span4Mux_v
    port map (
            O => \N__29068\,
            I => \N__29060\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29060\
        );

    \I__6619\ : Span4Mux_h
    port map (
            O => \N__29060\,
            I => \N__29057\
        );

    \I__6618\ : Odrv4
    port map (
            O => \N__29057\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_5\
        );

    \I__6617\ : InMux
    port map (
            O => \N__29054\,
            I => \N__29048\
        );

    \I__6616\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29048\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__29048\,
            I => \N__29045\
        );

    \I__6614\ : Span4Mux_s3_h
    port map (
            O => \N__29045\,
            I => \N__29042\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__29042\,
            I => \N__29039\
        );

    \I__6612\ : Odrv4
    port map (
            O => \N__29039\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_6\
        );

    \I__6611\ : CEMux
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__29033\,
            I => \N__29030\
        );

    \I__6609\ : Span4Mux_v
    port map (
            O => \N__29030\,
            I => \N__29027\
        );

    \I__6608\ : Span4Mux_h
    port map (
            O => \N__29027\,
            I => \N__29024\
        );

    \I__6607\ : Span4Mux_h
    port map (
            O => \N__29024\,
            I => \N__29021\
        );

    \I__6606\ : Odrv4
    port map (
            O => \N__29021\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe26\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__29018\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_7_cascade_\
        );

    \I__6604\ : InMux
    port map (
            O => \N__29015\,
            I => \N__29009\
        );

    \I__6603\ : InMux
    port map (
            O => \N__29014\,
            I => \N__29006\
        );

    \I__6602\ : InMux
    port map (
            O => \N__29013\,
            I => \N__28994\
        );

    \I__6601\ : InMux
    port map (
            O => \N__29012\,
            I => \N__28991\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__29009\,
            I => \N__28988\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__29006\,
            I => \N__28985\
        );

    \I__6598\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28982\
        );

    \I__6597\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28979\
        );

    \I__6596\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28975\
        );

    \I__6595\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28970\
        );

    \I__6594\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28965\
        );

    \I__6593\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28960\
        );

    \I__6592\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28960\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__28998\,
            I => \N__28951\
        );

    \I__6590\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28946\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__28994\,
            I => \N__28921\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28918\
        );

    \I__6587\ : Span4Mux_s1_h
    port map (
            O => \N__28988\,
            I => \N__28909\
        );

    \I__6586\ : Span4Mux_v
    port map (
            O => \N__28985\,
            I => \N__28909\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28909\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__28979\,
            I => \N__28909\
        );

    \I__6583\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28906\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__28975\,
            I => \N__28903\
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__28974\,
            I => \N__28900\
        );

    \I__6580\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28897\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__28970\,
            I => \N__28894\
        );

    \I__6578\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28890\
        );

    \I__6577\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28886\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__28965\,
            I => \N__28882\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__28960\,
            I => \N__28879\
        );

    \I__6574\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28870\
        );

    \I__6573\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28870\
        );

    \I__6572\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28870\
        );

    \I__6571\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28870\
        );

    \I__6570\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28867\
        );

    \I__6569\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28858\
        );

    \I__6568\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28858\
        );

    \I__6567\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28858\
        );

    \I__6566\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28858\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__28946\,
            I => \N__28855\
        );

    \I__6564\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28850\
        );

    \I__6563\ : InMux
    port map (
            O => \N__28944\,
            I => \N__28850\
        );

    \I__6562\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28841\
        );

    \I__6561\ : InMux
    port map (
            O => \N__28942\,
            I => \N__28841\
        );

    \I__6560\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28841\
        );

    \I__6559\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28841\
        );

    \I__6558\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28828\
        );

    \I__6557\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28828\
        );

    \I__6556\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28828\
        );

    \I__6555\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28828\
        );

    \I__6554\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28828\
        );

    \I__6553\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28828\
        );

    \I__6552\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28819\
        );

    \I__6551\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28819\
        );

    \I__6550\ : InMux
    port map (
            O => \N__28931\,
            I => \N__28819\
        );

    \I__6549\ : InMux
    port map (
            O => \N__28930\,
            I => \N__28819\
        );

    \I__6548\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28814\
        );

    \I__6547\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28814\
        );

    \I__6546\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28809\
        );

    \I__6545\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28809\
        );

    \I__6544\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28806\
        );

    \I__6543\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28803\
        );

    \I__6542\ : Span4Mux_s1_h
    port map (
            O => \N__28921\,
            I => \N__28794\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__28918\,
            I => \N__28794\
        );

    \I__6540\ : Span4Mux_v
    port map (
            O => \N__28909\,
            I => \N__28794\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__28906\,
            I => \N__28794\
        );

    \I__6538\ : Span4Mux_s2_h
    port map (
            O => \N__28903\,
            I => \N__28791\
        );

    \I__6537\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28788\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__28897\,
            I => \N__28785\
        );

    \I__6535\ : Span4Mux_v
    port map (
            O => \N__28894\,
            I => \N__28782\
        );

    \I__6534\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28775\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28771\
        );

    \I__6532\ : InMux
    port map (
            O => \N__28889\,
            I => \N__28768\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__28886\,
            I => \N__28763\
        );

    \I__6530\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28760\
        );

    \I__6529\ : Span4Mux_v
    port map (
            O => \N__28882\,
            I => \N__28749\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__28879\,
            I => \N__28749\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28749\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28749\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28749\
        );

    \I__6524\ : Span4Mux_h
    port map (
            O => \N__28855\,
            I => \N__28740\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__28850\,
            I => \N__28740\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28740\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28740\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28733\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28733\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28733\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__28806\,
            I => \N__28726\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28726\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__28794\,
            I => \N__28726\
        );

    \I__6514\ : Sp12to4
    port map (
            O => \N__28791\,
            I => \N__28723\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__28788\,
            I => \N__28716\
        );

    \I__6512\ : Span4Mux_v
    port map (
            O => \N__28785\,
            I => \N__28716\
        );

    \I__6511\ : Span4Mux_h
    port map (
            O => \N__28782\,
            I => \N__28716\
        );

    \I__6510\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28707\
        );

    \I__6509\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28707\
        );

    \I__6508\ : InMux
    port map (
            O => \N__28779\,
            I => \N__28707\
        );

    \I__6507\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28707\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__28775\,
            I => \N__28704\
        );

    \I__6505\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28701\
        );

    \I__6504\ : Span4Mux_v
    port map (
            O => \N__28771\,
            I => \N__28696\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28696\
        );

    \I__6502\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28691\
        );

    \I__6501\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28691\
        );

    \I__6500\ : Span4Mux_v
    port map (
            O => \N__28763\,
            I => \N__28684\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__28760\,
            I => \N__28684\
        );

    \I__6498\ : Span4Mux_v
    port map (
            O => \N__28749\,
            I => \N__28684\
        );

    \I__6497\ : Span4Mux_v
    port map (
            O => \N__28740\,
            I => \N__28677\
        );

    \I__6496\ : Span4Mux_h
    port map (
            O => \N__28733\,
            I => \N__28677\
        );

    \I__6495\ : Span4Mux_h
    port map (
            O => \N__28726\,
            I => \N__28677\
        );

    \I__6494\ : Odrv12
    port map (
            O => \N__28723\,
            I => instruction_5
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__28716\,
            I => instruction_5
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__28707\,
            I => instruction_5
        );

    \I__6491\ : Odrv4
    port map (
            O => \N__28704\,
            I => instruction_5
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__28701\,
            I => instruction_5
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__28696\,
            I => instruction_5
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__28691\,
            I => instruction_5
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__28684\,
            I => instruction_5
        );

    \I__6486\ : Odrv4
    port map (
            O => \N__28677\,
            I => instruction_5
        );

    \I__6485\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28642\
        );

    \I__6484\ : CascadeMux
    port map (
            O => \N__28657\,
            I => \N__28634\
        );

    \I__6483\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28628\
        );

    \I__6482\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28628\
        );

    \I__6481\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28623\
        );

    \I__6480\ : InMux
    port map (
            O => \N__28653\,
            I => \N__28623\
        );

    \I__6479\ : InMux
    port map (
            O => \N__28652\,
            I => \N__28608\
        );

    \I__6478\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28608\
        );

    \I__6477\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28603\
        );

    \I__6476\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28603\
        );

    \I__6475\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28593\
        );

    \I__6474\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28593\
        );

    \I__6473\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28588\
        );

    \I__6472\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28588\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__28642\,
            I => \N__28582\
        );

    \I__6470\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28577\
        );

    \I__6469\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28577\
        );

    \I__6468\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28572\
        );

    \I__6467\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28563\
        );

    \I__6466\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28563\
        );

    \I__6465\ : InMux
    port map (
            O => \N__28634\,
            I => \N__28563\
        );

    \I__6464\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28563\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__28628\,
            I => \N__28551\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__28623\,
            I => \N__28551\
        );

    \I__6461\ : InMux
    port map (
            O => \N__28622\,
            I => \N__28546\
        );

    \I__6460\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28546\
        );

    \I__6459\ : InMux
    port map (
            O => \N__28620\,
            I => \N__28539\
        );

    \I__6458\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28539\
        );

    \I__6457\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28534\
        );

    \I__6456\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28534\
        );

    \I__6455\ : InMux
    port map (
            O => \N__28616\,
            I => \N__28529\
        );

    \I__6454\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28529\
        );

    \I__6453\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28522\
        );

    \I__6452\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28522\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28519\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__28603\,
            I => \N__28516\
        );

    \I__6449\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28511\
        );

    \I__6448\ : InMux
    port map (
            O => \N__28601\,
            I => \N__28511\
        );

    \I__6447\ : InMux
    port map (
            O => \N__28600\,
            I => \N__28506\
        );

    \I__6446\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28506\
        );

    \I__6445\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28503\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__28593\,
            I => \N__28498\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__28588\,
            I => \N__28498\
        );

    \I__6442\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28495\
        );

    \I__6441\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28490\
        );

    \I__6440\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28490\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__28582\,
            I => \N__28485\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__28577\,
            I => \N__28485\
        );

    \I__6437\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28480\
        );

    \I__6436\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28480\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__28572\,
            I => \N__28475\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28475\
        );

    \I__6433\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28468\
        );

    \I__6432\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28468\
        );

    \I__6431\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28468\
        );

    \I__6430\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28461\
        );

    \I__6429\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28461\
        );

    \I__6428\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28461\
        );

    \I__6427\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28458\
        );

    \I__6426\ : Span4Mux_v
    port map (
            O => \N__28551\,
            I => \N__28453\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__28546\,
            I => \N__28453\
        );

    \I__6424\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28448\
        );

    \I__6423\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28448\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28443\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__28534\,
            I => \N__28443\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__28529\,
            I => \N__28437\
        );

    \I__6419\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28432\
        );

    \I__6418\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28432\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28429\
        );

    \I__6416\ : Span4Mux_v
    port map (
            O => \N__28519\,
            I => \N__28420\
        );

    \I__6415\ : Span4Mux_v
    port map (
            O => \N__28516\,
            I => \N__28420\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28415\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__28506\,
            I => \N__28415\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__28503\,
            I => \N__28406\
        );

    \I__6411\ : Span4Mux_v
    port map (
            O => \N__28498\,
            I => \N__28406\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__28495\,
            I => \N__28406\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28406\
        );

    \I__6408\ : Span4Mux_s3_h
    port map (
            O => \N__28485\,
            I => \N__28401\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__28480\,
            I => \N__28401\
        );

    \I__6406\ : Span4Mux_v
    port map (
            O => \N__28475\,
            I => \N__28392\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__28468\,
            I => \N__28392\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__28461\,
            I => \N__28392\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__28458\,
            I => \N__28392\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__28453\,
            I => \N__28385\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__28448\,
            I => \N__28385\
        );

    \I__6400\ : Span4Mux_v
    port map (
            O => \N__28443\,
            I => \N__28385\
        );

    \I__6399\ : InMux
    port map (
            O => \N__28442\,
            I => \N__28378\
        );

    \I__6398\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28378\
        );

    \I__6397\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28378\
        );

    \I__6396\ : Span4Mux_s1_h
    port map (
            O => \N__28437\,
            I => \N__28373\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__28432\,
            I => \N__28373\
        );

    \I__6394\ : Span4Mux_v
    port map (
            O => \N__28429\,
            I => \N__28370\
        );

    \I__6393\ : InMux
    port map (
            O => \N__28428\,
            I => \N__28365\
        );

    \I__6392\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28365\
        );

    \I__6391\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28360\
        );

    \I__6390\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28360\
        );

    \I__6389\ : Span4Mux_h
    port map (
            O => \N__28420\,
            I => \N__28353\
        );

    \I__6388\ : Span4Mux_v
    port map (
            O => \N__28415\,
            I => \N__28353\
        );

    \I__6387\ : Span4Mux_v
    port map (
            O => \N__28406\,
            I => \N__28353\
        );

    \I__6386\ : Span4Mux_v
    port map (
            O => \N__28401\,
            I => \N__28346\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__28392\,
            I => \N__28346\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__28385\,
            I => \N__28346\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__28378\,
            I => instruction_6
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__28373\,
            I => instruction_6
        );

    \I__6381\ : Odrv4
    port map (
            O => \N__28370\,
            I => instruction_6
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__28365\,
            I => instruction_6
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__28360\,
            I => instruction_6
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__28353\,
            I => instruction_6
        );

    \I__6377\ : Odrv4
    port map (
            O => \N__28346\,
            I => instruction_6
        );

    \I__6376\ : InMux
    port map (
            O => \N__28331\,
            I => \N__28328\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__6374\ : Span4Mux_s0_h
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__6373\ : Odrv4
    port map (
            O => \N__28322\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_7\
        );

    \I__6372\ : CascadeMux
    port map (
            O => \N__28319\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_7_cascade_\
        );

    \I__6371\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__28313\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_7\
        );

    \I__6369\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28307\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__28307\,
            I => \N__28304\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__28304\,
            I => \N__28301\
        );

    \I__6366\ : Span4Mux_h
    port map (
            O => \N__28301\,
            I => \N__28298\
        );

    \I__6365\ : Span4Mux_h
    port map (
            O => \N__28298\,
            I => \N__28295\
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__28295\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_7\
        );

    \I__6363\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28288\
        );

    \I__6362\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28285\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__28288\,
            I => \N__28280\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__28285\,
            I => \N__28280\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__28280\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_7\
        );

    \I__6358\ : CascadeMux
    port map (
            O => \N__28277\,
            I => \N__28274\
        );

    \I__6357\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28268\
        );

    \I__6356\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28268\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__6354\ : Odrv12
    port map (
            O => \N__28265\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_7\
        );

    \I__6353\ : CascadeMux
    port map (
            O => \N__28262\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_7_cascade_\
        );

    \I__6352\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28256\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__28256\,
            I => \N__28253\
        );

    \I__6350\ : Span4Mux_h
    port map (
            O => \N__28253\,
            I => \N__28250\
        );

    \I__6349\ : Span4Mux_h
    port map (
            O => \N__28250\,
            I => \N__28247\
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__28247\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI0NMM1_7\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__28244\,
            I => \N__28241\
        );

    \I__6346\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28237\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__28240\,
            I => \N__28234\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__28237\,
            I => \N__28231\
        );

    \I__6343\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28228\
        );

    \I__6342\ : Span4Mux_h
    port map (
            O => \N__28231\,
            I => \N__28225\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__28228\,
            I => \N__28222\
        );

    \I__6340\ : Odrv4
    port map (
            O => \N__28225\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4\
        );

    \I__6339\ : Odrv4
    port map (
            O => \N__28222\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__28217\,
            I => \N__28213\
        );

    \I__6337\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28208\
        );

    \I__6336\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28208\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__28208\,
            I => \N__28205\
        );

    \I__6334\ : Span4Mux_v
    port map (
            O => \N__28205\,
            I => \N__28202\
        );

    \I__6333\ : Odrv4
    port map (
            O => \N__28202\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_5\
        );

    \I__6332\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28195\
        );

    \I__6331\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28192\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__28195\,
            I => \N__28187\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__28192\,
            I => \N__28187\
        );

    \I__6328\ : Span4Mux_h
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__28184\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_6\
        );

    \I__6326\ : CEMux
    port map (
            O => \N__28181\,
            I => \N__28178\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__28178\,
            I => \N__28175\
        );

    \I__6324\ : Span4Mux_s3_h
    port map (
            O => \N__28175\,
            I => \N__28172\
        );

    \I__6323\ : Span4Mux_v
    port map (
            O => \N__28172\,
            I => \N__28169\
        );

    \I__6322\ : Span4Mux_h
    port map (
            O => \N__28169\,
            I => \N__28166\
        );

    \I__6321\ : Odrv4
    port map (
            O => \N__28166\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe25\
        );

    \I__6320\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28160\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__28160\,
            I => \N__28156\
        );

    \I__6318\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28153\
        );

    \I__6317\ : Span4Mux_h
    port map (
            O => \N__28156\,
            I => \N__28150\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__28153\,
            I => \N__28147\
        );

    \I__6315\ : Odrv4
    port map (
            O => \N__28150\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0\
        );

    \I__6314\ : Odrv12
    port map (
            O => \N__28147\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0\
        );

    \I__6313\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28136\
        );

    \I__6312\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28136\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__28136\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_1\
        );

    \I__6310\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28130\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__28130\,
            I => \N__28126\
        );

    \I__6308\ : CascadeMux
    port map (
            O => \N__28129\,
            I => \N__28123\
        );

    \I__6307\ : Span4Mux_v
    port map (
            O => \N__28126\,
            I => \N__28120\
        );

    \I__6306\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28117\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__28120\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__28117\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2\
        );

    \I__6303\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28109\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__28109\,
            I => \N__28105\
        );

    \I__6301\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28102\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__28105\,
            I => \N__28099\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28096\
        );

    \I__6298\ : Odrv4
    port map (
            O => \N__28099\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__28096\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3\
        );

    \I__6296\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28088\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__28088\,
            I => \N__28085\
        );

    \I__6294\ : Span4Mux_v
    port map (
            O => \N__28085\,
            I => \N__28081\
        );

    \I__6293\ : InMux
    port map (
            O => \N__28084\,
            I => \N__28078\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__28081\,
            I => \N__28075\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__28078\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4\
        );

    \I__6290\ : Odrv4
    port map (
            O => \N__28075\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4\
        );

    \I__6289\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28064\
        );

    \I__6288\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28064\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__28064\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_3\
        );

    \I__6286\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28057\
        );

    \I__6285\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28054\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28051\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__28054\,
            I => \N__28048\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__28051\,
            I => \N__28045\
        );

    \I__6281\ : Span4Mux_v
    port map (
            O => \N__28048\,
            I => \N__28042\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__28045\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__28042\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4\
        );

    \I__6278\ : InMux
    port map (
            O => \N__28037\,
            I => \N__28031\
        );

    \I__6277\ : InMux
    port map (
            O => \N__28036\,
            I => \N__28031\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__28031\,
            I => \N__28028\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__28028\,
            I => \N__28025\
        );

    \I__6274\ : Odrv4
    port map (
            O => \N__28025\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_5\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__28022\,
            I => \N__28019\
        );

    \I__6272\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28013\
        );

    \I__6271\ : InMux
    port map (
            O => \N__28018\,
            I => \N__28013\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__6269\ : Span4Mux_h
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__28007\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_6\
        );

    \I__6267\ : CEMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__28001\,
            I => \N__27998\
        );

    \I__6265\ : Span4Mux_s0_h
    port map (
            O => \N__27998\,
            I => \N__27995\
        );

    \I__6264\ : Span4Mux_h
    port map (
            O => \N__27995\,
            I => \N__27992\
        );

    \I__6263\ : Odrv4
    port map (
            O => \N__27992\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe24\
        );

    \I__6262\ : CascadeMux
    port map (
            O => \N__27989\,
            I => \N__27985\
        );

    \I__6261\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27980\
        );

    \I__6260\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27980\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__27980\,
            I => \N__27977\
        );

    \I__6258\ : Span4Mux_h
    port map (
            O => \N__27977\,
            I => \N__27974\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__27974\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_0\
        );

    \I__6256\ : CascadeMux
    port map (
            O => \N__27971\,
            I => \N__27968\
        );

    \I__6255\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27964\
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__27967\,
            I => \N__27961\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__27964\,
            I => \N__27958\
        );

    \I__6252\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27955\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__27958\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__27955\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1\
        );

    \I__6249\ : InMux
    port map (
            O => \N__27950\,
            I => \N__27944\
        );

    \I__6248\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27944\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__27944\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_2\
        );

    \I__6246\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27935\
        );

    \I__6245\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27935\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__27935\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_3\
        );

    \I__6243\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27929\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27925\
        );

    \I__6241\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27922\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__27925\,
            I => \N__27917\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__27922\,
            I => \N__27917\
        );

    \I__6238\ : Span4Mux_v
    port map (
            O => \N__27917\,
            I => \N__27914\
        );

    \I__6237\ : Odrv4
    port map (
            O => \N__27914\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_3\
        );

    \I__6236\ : CascadeMux
    port map (
            O => \N__27911\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_3_cascade_\
        );

    \I__6235\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27904\
        );

    \I__6234\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27901\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__27904\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__27901\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3\
        );

    \I__6231\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__27893\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIKIUU1_3\
        );

    \I__6229\ : CascadeMux
    port map (
            O => \N__27890\,
            I => \N__27887\
        );

    \I__6228\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27883\
        );

    \I__6227\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27880\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__27883\,
            I => \N__27877\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__27880\,
            I => \N__27874\
        );

    \I__6224\ : Span4Mux_v
    port map (
            O => \N__27877\,
            I => \N__27869\
        );

    \I__6223\ : Span4Mux_v
    port map (
            O => \N__27874\,
            I => \N__27869\
        );

    \I__6222\ : Odrv4
    port map (
            O => \N__27869\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_3\
        );

    \I__6221\ : InMux
    port map (
            O => \N__27866\,
            I => \N__27862\
        );

    \I__6220\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27859\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__27862\,
            I => \N__27856\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__27859\,
            I => \N__27853\
        );

    \I__6217\ : Span4Mux_s3_h
    port map (
            O => \N__27856\,
            I => \N__27850\
        );

    \I__6216\ : Span4Mux_s2_h
    port map (
            O => \N__27853\,
            I => \N__27847\
        );

    \I__6215\ : Odrv4
    port map (
            O => \N__27850\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__27847\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3\
        );

    \I__6213\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27839\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__27839\,
            I => \N__27836\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__27836\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_3\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__27833\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_3_cascade_\
        );

    \I__6209\ : CascadeMux
    port map (
            O => \N__27830\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_3_cascade_\
        );

    \I__6208\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27824\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__27824\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_3\
        );

    \I__6206\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27818\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__6204\ : Span4Mux_h
    port map (
            O => \N__27815\,
            I => \N__27812\
        );

    \I__6203\ : Odrv4
    port map (
            O => \N__27812\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_3\
        );

    \I__6202\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27805\
        );

    \I__6201\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27802\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__27805\,
            I => \N__27799\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__27802\,
            I => \N__27796\
        );

    \I__6198\ : Span12Mux_s1_h
    port map (
            O => \N__27799\,
            I => \N__27791\
        );

    \I__6197\ : Span12Mux_s7_v
    port map (
            O => \N__27796\,
            I => \N__27791\
        );

    \I__6196\ : Odrv12
    port map (
            O => \N__27791\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_2\
        );

    \I__6195\ : CEMux
    port map (
            O => \N__27788\,
            I => \N__27785\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__27785\,
            I => \N__27782\
        );

    \I__6193\ : Span4Mux_v
    port map (
            O => \N__27782\,
            I => \N__27778\
        );

    \I__6192\ : CEMux
    port map (
            O => \N__27781\,
            I => \N__27775\
        );

    \I__6191\ : Span4Mux_h
    port map (
            O => \N__27778\,
            I => \N__27771\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__27775\,
            I => \N__27768\
        );

    \I__6189\ : CEMux
    port map (
            O => \N__27774\,
            I => \N__27765\
        );

    \I__6188\ : Span4Mux_v
    port map (
            O => \N__27771\,
            I => \N__27762\
        );

    \I__6187\ : Span4Mux_h
    port map (
            O => \N__27768\,
            I => \N__27759\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__27765\,
            I => \N__27756\
        );

    \I__6185\ : Odrv4
    port map (
            O => \N__27762\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31\
        );

    \I__6184\ : Odrv4
    port map (
            O => \N__27759\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31\
        );

    \I__6183\ : Odrv12
    port map (
            O => \N__27756\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31\
        );

    \I__6182\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27743\
        );

    \I__6181\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27743\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__27743\,
            I => \N__27740\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__27740\,
            I => \N__27737\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__27737\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_0\
        );

    \I__6177\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27731\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__27731\,
            I => \N__27728\
        );

    \I__6175\ : Span4Mux_v
    port map (
            O => \N__27728\,
            I => \N__27724\
        );

    \I__6174\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27721\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__27724\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__27721\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1\
        );

    \I__6171\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27710\
        );

    \I__6170\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27710\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__27710\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_2\
        );

    \I__6168\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27703\
        );

    \I__6167\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27700\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__27703\,
            I => \N__27697\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__27700\,
            I => \N__27692\
        );

    \I__6164\ : Span4Mux_h
    port map (
            O => \N__27697\,
            I => \N__27692\
        );

    \I__6163\ : Span4Mux_h
    port map (
            O => \N__27692\,
            I => \N__27689\
        );

    \I__6162\ : Odrv4
    port map (
            O => \N__27689\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_4\
        );

    \I__6161\ : CEMux
    port map (
            O => \N__27686\,
            I => \N__27683\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__27683\,
            I => \N__27680\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__27680\,
            I => \N__27676\
        );

    \I__6158\ : CEMux
    port map (
            O => \N__27679\,
            I => \N__27673\
        );

    \I__6157\ : Span4Mux_s0_h
    port map (
            O => \N__27676\,
            I => \N__27670\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__27673\,
            I => \N__27667\
        );

    \I__6155\ : Span4Mux_h
    port map (
            O => \N__27670\,
            I => \N__27664\
        );

    \I__6154\ : Span4Mux_s1_v
    port map (
            O => \N__27667\,
            I => \N__27661\
        );

    \I__6153\ : Span4Mux_h
    port map (
            O => \N__27664\,
            I => \N__27658\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__27661\,
            I => \N__27655\
        );

    \I__6151\ : Span4Mux_s3_h
    port map (
            O => \N__27658\,
            I => \N__27652\
        );

    \I__6150\ : Odrv4
    port map (
            O => \N__27655\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18\
        );

    \I__6149\ : Odrv4
    port map (
            O => \N__27652\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__27647\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_3_cascade_\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__27644\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI06K32_3_cascade_\
        );

    \I__6146\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27637\
        );

    \I__6145\ : InMux
    port map (
            O => \N__27640\,
            I => \N__27633\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__27637\,
            I => \N__27625\
        );

    \I__6143\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27621\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__27633\,
            I => \N__27618\
        );

    \I__6141\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27615\
        );

    \I__6140\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27612\
        );

    \I__6139\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27606\
        );

    \I__6138\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27602\
        );

    \I__6137\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27599\
        );

    \I__6136\ : Span4Mux_v
    port map (
            O => \N__27625\,
            I => \N__27596\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__27624\,
            I => \N__27591\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27587\
        );

    \I__6133\ : Span4Mux_v
    port map (
            O => \N__27618\,
            I => \N__27582\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__27615\,
            I => \N__27582\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__27612\,
            I => \N__27579\
        );

    \I__6130\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27574\
        );

    \I__6129\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27574\
        );

    \I__6128\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27571\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__27606\,
            I => \N__27568\
        );

    \I__6126\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27565\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__27602\,
            I => \N__27559\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__27599\,
            I => \N__27559\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__27596\,
            I => \N__27556\
        );

    \I__6122\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27551\
        );

    \I__6121\ : InMux
    port map (
            O => \N__27594\,
            I => \N__27551\
        );

    \I__6120\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27545\
        );

    \I__6119\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27545\
        );

    \I__6118\ : Span4Mux_s2_h
    port map (
            O => \N__27587\,
            I => \N__27542\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__27582\,
            I => \N__27536\
        );

    \I__6116\ : Span4Mux_h
    port map (
            O => \N__27579\,
            I => \N__27533\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27524\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__27571\,
            I => \N__27524\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__27568\,
            I => \N__27524\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27524\
        );

    \I__6111\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27521\
        );

    \I__6110\ : Span4Mux_h
    port map (
            O => \N__27559\,
            I => \N__27518\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__27556\,
            I => \N__27513\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__27551\,
            I => \N__27513\
        );

    \I__6107\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27510\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27505\
        );

    \I__6105\ : Span4Mux_h
    port map (
            O => \N__27542\,
            I => \N__27505\
        );

    \I__6104\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27502\
        );

    \I__6103\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27499\
        );

    \I__6102\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27496\
        );

    \I__6101\ : Span4Mux_v
    port map (
            O => \N__27536\,
            I => \N__27493\
        );

    \I__6100\ : Span4Mux_v
    port map (
            O => \N__27533\,
            I => \N__27486\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__27524\,
            I => \N__27486\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27486\
        );

    \I__6097\ : Span4Mux_v
    port map (
            O => \N__27518\,
            I => \N__27479\
        );

    \I__6096\ : Span4Mux_h
    port map (
            O => \N__27513\,
            I => \N__27479\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__27510\,
            I => \N__27479\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__27505\,
            I => \N__27472\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__27502\,
            I => \N__27472\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__27499\,
            I => \N__27472\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__27496\,
            I => instruction_10
        );

    \I__6090\ : Odrv4
    port map (
            O => \N__27493\,
            I => instruction_10
        );

    \I__6089\ : Odrv4
    port map (
            O => \N__27486\,
            I => instruction_10
        );

    \I__6088\ : Odrv4
    port map (
            O => \N__27479\,
            I => instruction_10
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__27472\,
            I => instruction_10
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__27461\,
            I => \N__27457\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__27460\,
            I => \N__27436\
        );

    \I__6084\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27425\
        );

    \I__6083\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27410\
        );

    \I__6082\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27410\
        );

    \I__6081\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27410\
        );

    \I__6080\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27410\
        );

    \I__6079\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27410\
        );

    \I__6078\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27410\
        );

    \I__6077\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27410\
        );

    \I__6076\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27395\
        );

    \I__6075\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27395\
        );

    \I__6074\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27395\
        );

    \I__6073\ : InMux
    port map (
            O => \N__27446\,
            I => \N__27395\
        );

    \I__6072\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27395\
        );

    \I__6071\ : InMux
    port map (
            O => \N__27444\,
            I => \N__27395\
        );

    \I__6070\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27395\
        );

    \I__6069\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27381\
        );

    \I__6068\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27374\
        );

    \I__6067\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27374\
        );

    \I__6066\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27374\
        );

    \I__6065\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27371\
        );

    \I__6064\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27354\
        );

    \I__6063\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27354\
        );

    \I__6062\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27354\
        );

    \I__6061\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27354\
        );

    \I__6060\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27354\
        );

    \I__6059\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27354\
        );

    \I__6058\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27354\
        );

    \I__6057\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27354\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__27425\,
            I => \N__27347\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__27410\,
            I => \N__27347\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27347\
        );

    \I__6053\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27332\
        );

    \I__6052\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27332\
        );

    \I__6051\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27332\
        );

    \I__6050\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27332\
        );

    \I__6049\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27332\
        );

    \I__6048\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27332\
        );

    \I__6047\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27332\
        );

    \I__6046\ : InMux
    port map (
            O => \N__27387\,
            I => \N__27327\
        );

    \I__6045\ : InMux
    port map (
            O => \N__27386\,
            I => \N__27327\
        );

    \I__6044\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27322\
        );

    \I__6043\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27322\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__27381\,
            I => \N__27317\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__27374\,
            I => \N__27309\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__27371\,
            I => \N__27298\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__27354\,
            I => \N__27298\
        );

    \I__6038\ : Span4Mux_v
    port map (
            O => \N__27347\,
            I => \N__27298\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__27332\,
            I => \N__27298\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__27327\,
            I => \N__27298\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27295\
        );

    \I__6034\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27290\
        );

    \I__6033\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27290\
        );

    \I__6032\ : Span4Mux_v
    port map (
            O => \N__27317\,
            I => \N__27282\
        );

    \I__6031\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27279\
        );

    \I__6030\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27268\
        );

    \I__6029\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27268\
        );

    \I__6028\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27263\
        );

    \I__6027\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27263\
        );

    \I__6026\ : Span4Mux_h
    port map (
            O => \N__27309\,
            I => \N__27260\
        );

    \I__6025\ : Span4Mux_h
    port map (
            O => \N__27298\,
            I => \N__27253\
        );

    \I__6024\ : Span4Mux_s3_v
    port map (
            O => \N__27295\,
            I => \N__27253\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__27290\,
            I => \N__27253\
        );

    \I__6022\ : InMux
    port map (
            O => \N__27289\,
            I => \N__27248\
        );

    \I__6021\ : InMux
    port map (
            O => \N__27288\,
            I => \N__27245\
        );

    \I__6020\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27242\
        );

    \I__6019\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27239\
        );

    \I__6018\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27236\
        );

    \I__6017\ : Span4Mux_s1_h
    port map (
            O => \N__27282\,
            I => \N__27231\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__27279\,
            I => \N__27231\
        );

    \I__6015\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27226\
        );

    \I__6014\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27226\
        );

    \I__6013\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27217\
        );

    \I__6012\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27217\
        );

    \I__6011\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27217\
        );

    \I__6010\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27217\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__27268\,
            I => \N__27212\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27212\
        );

    \I__6007\ : Span4Mux_h
    port map (
            O => \N__27260\,
            I => \N__27207\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__27253\,
            I => \N__27207\
        );

    \I__6005\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27200\
        );

    \I__6004\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27200\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__27248\,
            I => \N__27193\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__27245\,
            I => \N__27193\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27193\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__27239\,
            I => \N__27188\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__27236\,
            I => \N__27183\
        );

    \I__5998\ : Span4Mux_h
    port map (
            O => \N__27231\,
            I => \N__27178\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27226\,
            I => \N__27178\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__27217\,
            I => \N__27173\
        );

    \I__5995\ : Span4Mux_v
    port map (
            O => \N__27212\,
            I => \N__27173\
        );

    \I__5994\ : IoSpan4Mux
    port map (
            O => \N__27207\,
            I => \N__27170\
        );

    \I__5993\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27165\
        );

    \I__5992\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27165\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__27200\,
            I => \N__27160\
        );

    \I__5990\ : Span4Mux_v
    port map (
            O => \N__27193\,
            I => \N__27160\
        );

    \I__5989\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27155\
        );

    \I__5988\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27155\
        );

    \I__5987\ : Span12Mux_s9_h
    port map (
            O => \N__27188\,
            I => \N__27152\
        );

    \I__5986\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27147\
        );

    \I__5985\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27147\
        );

    \I__5984\ : Span4Mux_h
    port map (
            O => \N__27183\,
            I => \N__27142\
        );

    \I__5983\ : Span4Mux_h
    port map (
            O => \N__27178\,
            I => \N__27142\
        );

    \I__5982\ : Span4Mux_h
    port map (
            O => \N__27173\,
            I => \N__27131\
        );

    \I__5981\ : Span4Mux_s1_h
    port map (
            O => \N__27170\,
            I => \N__27131\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__27165\,
            I => \N__27131\
        );

    \I__5979\ : Span4Mux_h
    port map (
            O => \N__27160\,
            I => \N__27131\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__27155\,
            I => \N__27131\
        );

    \I__5977\ : Odrv12
    port map (
            O => \N__27152\,
            I => instruction_11
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__27147\,
            I => instruction_11
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__27142\,
            I => instruction_11
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__27131\,
            I => instruction_11
        );

    \I__5973\ : InMux
    port map (
            O => \N__27122\,
            I => \N__27119\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__5971\ : Odrv12
    port map (
            O => \N__27116\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIE0IQ1_3\
        );

    \I__5970\ : CascadeMux
    port map (
            O => \N__27113\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_3_cascade_\
        );

    \I__5969\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27104\
        );

    \I__5967\ : Span4Mux_v
    port map (
            O => \N__27104\,
            I => \N__27101\
        );

    \I__5966\ : Span4Mux_h
    port map (
            O => \N__27101\,
            I => \N__27098\
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__27098\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV1BI8_3\
        );

    \I__5964\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27091\
        );

    \I__5963\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27088\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__27091\,
            I => \N__27085\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__27088\,
            I => \N__27082\
        );

    \I__5960\ : Odrv12
    port map (
            O => \N__27085\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3\
        );

    \I__5959\ : Odrv4
    port map (
            O => \N__27082\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3\
        );

    \I__5958\ : CascadeMux
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__5957\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27071\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__27071\,
            I => \N__27068\
        );

    \I__5955\ : Odrv12
    port map (
            O => \N__27068\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_3\
        );

    \I__5954\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27062\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__27062\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIG6MM1_3\
        );

    \I__5952\ : InMux
    port map (
            O => \N__27059\,
            I => \N__27056\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__27056\,
            I => \N__27053\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__27053\,
            I => \N__27050\
        );

    \I__5949\ : Span4Mux_s0_h
    port map (
            O => \N__27050\,
            I => \N__27047\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__27047\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIASHQ1_2\
        );

    \I__5947\ : CascadeMux
    port map (
            O => \N__27044\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIC2MM1_2_cascade_\
        );

    \I__5946\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27035\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__5942\ : Odrv4
    port map (
            O => \N__27029\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFHAI8_2\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__5940\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27020\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__27020\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_2\
        );

    \I__5938\ : InMux
    port map (
            O => \N__27017\,
            I => \N__27014\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__27014\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIS1K32_2\
        );

    \I__5936\ : CascadeMux
    port map (
            O => \N__27011\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIGEUU1_2_cascade_\
        );

    \I__5935\ : InMux
    port map (
            O => \N__27008\,
            I => \N__27005\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__27005\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_2\
        );

    \I__5933\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26998\
        );

    \I__5932\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26995\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26992\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__26995\,
            I => \N__26989\
        );

    \I__5929\ : Span4Mux_h
    port map (
            O => \N__26992\,
            I => \N__26986\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__26989\,
            I => \N__26983\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__26986\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0\
        );

    \I__5926\ : Odrv4
    port map (
            O => \N__26983\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0\
        );

    \I__5925\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26974\
        );

    \I__5924\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26971\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__26974\,
            I => \N__26966\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__26971\,
            I => \N__26966\
        );

    \I__5921\ : Span4Mux_v
    port map (
            O => \N__26966\,
            I => \N__26963\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__26963\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_1\
        );

    \I__5919\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__26957\,
            I => \N__26953\
        );

    \I__5917\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26950\
        );

    \I__5916\ : Odrv4
    port map (
            O => \N__26953\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__26950\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__26945\,
            I => \N__26942\
        );

    \I__5913\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26939\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__26939\,
            I => \N__26936\
        );

    \I__5911\ : Odrv4
    port map (
            O => \N__26936\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_1\
        );

    \I__5910\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26929\
        );

    \I__5909\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26926\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__26929\,
            I => \N__26921\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__26926\,
            I => \N__26921\
        );

    \I__5906\ : Span4Mux_v
    port map (
            O => \N__26921\,
            I => \N__26918\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__26918\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_2\
        );

    \I__5904\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26911\
        );

    \I__5903\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26908\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__26911\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__26908\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2\
        );

    \I__5900\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26900\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__26900\,
            I => \N__26897\
        );

    \I__5898\ : Span4Mux_h
    port map (
            O => \N__26897\,
            I => \N__26894\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__26894\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_2\
        );

    \I__5896\ : InMux
    port map (
            O => \N__26891\,
            I => \N__26888\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__26888\,
            I => \N__26885\
        );

    \I__5894\ : IoSpan4Mux
    port map (
            O => \N__26885\,
            I => \N__26882\
        );

    \I__5893\ : Span4Mux_s3_h
    port map (
            O => \N__26882\,
            I => \N__26878\
        );

    \I__5892\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26875\
        );

    \I__5891\ : Sp12to4
    port map (
            O => \N__26878\,
            I => \N__26870\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__26875\,
            I => \N__26870\
        );

    \I__5889\ : Odrv12
    port map (
            O => \N__26870\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_1\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26867\,
            I => \N__26864\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__26864\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_1\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__26861\,
            I => \N__26857\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__5884\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26851\
        );

    \I__5883\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26848\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__26851\,
            I => \N__26845\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__26848\,
            I => \N__26842\
        );

    \I__5880\ : Span4Mux_v
    port map (
            O => \N__26845\,
            I => \N__26839\
        );

    \I__5879\ : Span4Mux_v
    port map (
            O => \N__26842\,
            I => \N__26836\
        );

    \I__5878\ : Span4Mux_v
    port map (
            O => \N__26839\,
            I => \N__26833\
        );

    \I__5877\ : Span4Mux_h
    port map (
            O => \N__26836\,
            I => \N__26830\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__26833\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1\
        );

    \I__5875\ : Odrv4
    port map (
            O => \N__26830\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1\
        );

    \I__5874\ : InMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__26822\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_295\
        );

    \I__5872\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__26816\,
            I => \N__26813\
        );

    \I__5870\ : Span4Mux_v
    port map (
            O => \N__26813\,
            I => \N__26809\
        );

    \I__5869\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26806\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__26809\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__26806\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__26801\,
            I => \N__26798\
        );

    \I__5865\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26795\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__26795\,
            I => \N__26791\
        );

    \I__5863\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26788\
        );

    \I__5862\ : Odrv4
    port map (
            O => \N__26791\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__26788\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__26783\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_1_cascade_\
        );

    \I__5859\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__26777\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_215\
        );

    \I__5857\ : InMux
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__26771\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_1\
        );

    \I__5855\ : CascadeMux
    port map (
            O => \N__26768\,
            I => \N__26765\
        );

    \I__5854\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__26762\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_239\
        );

    \I__5852\ : CascadeMux
    port map (
            O => \N__26759\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_2_cascade_\
        );

    \I__5851\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26753\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__26753\,
            I => \N__26749\
        );

    \I__5849\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26746\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__26749\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__26746\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2\
        );

    \I__5846\ : CascadeMux
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__5845\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26735\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26732\
        );

    \I__5843\ : Span4Mux_s2_h
    port map (
            O => \N__26732\,
            I => \N__26728\
        );

    \I__5842\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26725\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__26728\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__26725\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2\
        );

    \I__5839\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26713\
        );

    \I__5837\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26710\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__26713\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__26710\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__26705\,
            I => \N__26702\
        );

    \I__5833\ : InMux
    port map (
            O => \N__26702\,
            I => \N__26699\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26696\
        );

    \I__5831\ : Span4Mux_v
    port map (
            O => \N__26696\,
            I => \N__26693\
        );

    \I__5830\ : Odrv4
    port map (
            O => \N__26693\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_2\
        );

    \I__5829\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26686\
        );

    \I__5828\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26683\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__26686\,
            I => \N__26680\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__26683\,
            I => \N__26677\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__26680\,
            I => \N__26674\
        );

    \I__5824\ : Odrv12
    port map (
            O => \N__26677\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__26674\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__26669\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_4_cascade_\
        );

    \I__5821\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26663\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__26663\,
            I => \N__26660\
        );

    \I__5819\ : Span4Mux_v
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__5818\ : Span4Mux_h
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__26654\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIKAMM1_4\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__26651\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_1_cascade_\
        );

    \I__5815\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26644\
        );

    \I__5814\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26641\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__26644\,
            I => \N__26638\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__26641\,
            I => \N__26635\
        );

    \I__5811\ : Span4Mux_v
    port map (
            O => \N__26638\,
            I => \N__26632\
        );

    \I__5810\ : Span12Mux_s3_h
    port map (
            O => \N__26635\,
            I => \N__26629\
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__26632\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2\
        );

    \I__5808\ : Odrv12
    port map (
            O => \N__26629\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__26624\,
            I => \N__26621\
        );

    \I__5806\ : InMux
    port map (
            O => \N__26621\,
            I => \N__26617\
        );

    \I__5805\ : InMux
    port map (
            O => \N__26620\,
            I => \N__26614\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__26617\,
            I => \N__26609\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__26614\,
            I => \N__26609\
        );

    \I__5802\ : Odrv12
    port map (
            O => \N__26609\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_2\
        );

    \I__5801\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_2_cascade_\
        );

    \I__5800\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26599\
        );

    \I__5799\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26596\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__26599\,
            I => \N__26593\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26590\
        );

    \I__5796\ : Span4Mux_s2_h
    port map (
            O => \N__26593\,
            I => \N__26587\
        );

    \I__5795\ : Span4Mux_s2_h
    port map (
            O => \N__26590\,
            I => \N__26584\
        );

    \I__5794\ : Odrv4
    port map (
            O => \N__26587\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__26584\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2\
        );

    \I__5792\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26575\
        );

    \I__5791\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26572\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__26575\,
            I => \N__26569\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__26572\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1\
        );

    \I__5788\ : Odrv12
    port map (
            O => \N__26569\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1\
        );

    \I__5787\ : CascadeMux
    port map (
            O => \N__26564\,
            I => \N__26561\
        );

    \I__5786\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__26558\,
            I => \N__26555\
        );

    \I__5784\ : Odrv12
    port map (
            O => \N__26555\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_1\
        );

    \I__5783\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26549\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__5781\ : Span4Mux_h
    port map (
            O => \N__26546\,
            I => \N__26543\
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__26543\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1\
        );

    \I__5779\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26533\
        );

    \I__5777\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26530\
        );

    \I__5776\ : Span4Mux_v
    port map (
            O => \N__26533\,
            I => \N__26527\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__26530\,
            I => \N__26524\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__26527\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1\
        );

    \I__5773\ : Odrv12
    port map (
            O => \N__26524\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__26519\,
            I => \N__26516\
        );

    \I__5771\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26512\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__26515\,
            I => \N__26509\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__26512\,
            I => \N__26506\
        );

    \I__5768\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26503\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__26506\,
            I => \N__26500\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26497\
        );

    \I__5765\ : Span4Mux_v
    port map (
            O => \N__26500\,
            I => \N__26494\
        );

    \I__5764\ : Odrv12
    port map (
            O => \N__26497\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__26494\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1\
        );

    \I__5762\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26486\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26483\
        );

    \I__5760\ : Odrv12
    port map (
            O => \N__26483\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_271\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__26480\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_1_cascade_\
        );

    \I__5758\ : InMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__26474\,
            I => \N__26471\
        );

    \I__5756\ : Span4Mux_h
    port map (
            O => \N__26471\,
            I => \N__26468\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__26465\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_311\
        );

    \I__5753\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__26459\,
            I => \N__26455\
        );

    \I__5751\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26452\
        );

    \I__5750\ : Span4Mux_v
    port map (
            O => \N__26455\,
            I => \N__26447\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26447\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__26447\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_0\
        );

    \I__5747\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26440\
        );

    \I__5746\ : InMux
    port map (
            O => \N__26443\,
            I => \N__26437\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__26440\,
            I => \N__26434\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__26437\,
            I => \N__26431\
        );

    \I__5743\ : Span4Mux_h
    port map (
            O => \N__26434\,
            I => \N__26428\
        );

    \I__5742\ : Span4Mux_h
    port map (
            O => \N__26431\,
            I => \N__26425\
        );

    \I__5741\ : Odrv4
    port map (
            O => \N__26428\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__26425\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5\
        );

    \I__5739\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26414\
        );

    \I__5738\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26414\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__26414\,
            I => \N__26411\
        );

    \I__5736\ : Span12Mux_s6_v
    port map (
            O => \N__26411\,
            I => \N__26408\
        );

    \I__5735\ : Odrv12
    port map (
            O => \N__26408\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_6\
        );

    \I__5734\ : CEMux
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__5732\ : Span4Mux_v
    port map (
            O => \N__26399\,
            I => \N__26396\
        );

    \I__5731\ : Span4Mux_h
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__26393\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe27\
        );

    \I__5729\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__5727\ : Span4Mux_s3_h
    port map (
            O => \N__26384\,
            I => \N__26380\
        );

    \I__5726\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26377\
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__26380\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__26377\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__26372\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_3_cascade_\
        );

    \I__5722\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__26366\,
            I => \N__26362\
        );

    \I__5720\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26359\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__26362\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__26359\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__26354\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_2_cascade_\
        );

    \I__5716\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__26348\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_2\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__26345\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_2_cascade_\
        );

    \I__5713\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26336\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__5710\ : Span4Mux_v
    port map (
            O => \N__26333\,
            I => \N__26330\
        );

    \I__5709\ : Odrv4
    port map (
            O => \N__26330\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_2\
        );

    \I__5708\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__26324\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_2\
        );

    \I__5706\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__26318\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_2\
        );

    \I__5704\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26311\
        );

    \I__5703\ : InMux
    port map (
            O => \N__26314\,
            I => \N__26308\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__26311\,
            I => \N__26305\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__26308\,
            I => \N__26302\
        );

    \I__5700\ : Span4Mux_h
    port map (
            O => \N__26305\,
            I => \N__26297\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__26302\,
            I => \N__26297\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__26297\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_6\
        );

    \I__5697\ : CEMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__5695\ : Sp12to4
    port map (
            O => \N__26288\,
            I => \N__26285\
        );

    \I__5694\ : Odrv12
    port map (
            O => \N__26285\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe29\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__26282\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_3_cascade_\
        );

    \I__5692\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__5690\ : Odrv4
    port map (
            O => \N__26273\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_3\
        );

    \I__5689\ : CascadeMux
    port map (
            O => \N__26270\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_3_cascade_\
        );

    \I__5688\ : CascadeMux
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__5687\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__26252\,
            I => \N__26249\
        );

    \I__5682\ : Odrv4
    port map (
            O => \N__26249\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_3\
        );

    \I__5681\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26243\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__26243\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_3\
        );

    \I__5679\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26237\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__26237\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_3\
        );

    \I__5677\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26228\
        );

    \I__5676\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26228\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__26228\,
            I => \N__26225\
        );

    \I__5674\ : Span4Mux_s2_h
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__26222\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_3\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__26219\,
            I => \N__26216\
        );

    \I__5671\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26210\
        );

    \I__5670\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26210\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__26210\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_3\
        );

    \I__5668\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26204\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__26204\,
            I => \N__26201\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__26201\,
            I => \N__26197\
        );

    \I__5665\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26194\
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__26197\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__26194\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3\
        );

    \I__5662\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26186\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__26186\,
            I => \N__26182\
        );

    \I__5660\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26179\
        );

    \I__5659\ : Span4Mux_v
    port map (
            O => \N__26182\,
            I => \N__26176\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__26179\,
            I => \N__26173\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__26176\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__26173\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4\
        );

    \I__5655\ : CEMux
    port map (
            O => \N__26168\,
            I => \N__26164\
        );

    \I__5654\ : CEMux
    port map (
            O => \N__26167\,
            I => \N__26161\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__26164\,
            I => \N__26157\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__26161\,
            I => \N__26154\
        );

    \I__5651\ : CEMux
    port map (
            O => \N__26160\,
            I => \N__26151\
        );

    \I__5650\ : Sp12to4
    port map (
            O => \N__26157\,
            I => \N__26148\
        );

    \I__5649\ : Span4Mux_s3_v
    port map (
            O => \N__26154\,
            I => \N__26145\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__26151\,
            I => \N__26142\
        );

    \I__5647\ : Span12Mux_s5_h
    port map (
            O => \N__26148\,
            I => \N__26139\
        );

    \I__5646\ : Span4Mux_h
    port map (
            O => \N__26145\,
            I => \N__26136\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__26142\,
            I => \N__26133\
        );

    \I__5644\ : Odrv12
    port map (
            O => \N__26139\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3\
        );

    \I__5643\ : Odrv4
    port map (
            O => \N__26136\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__26133\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3\
        );

    \I__5641\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26122\
        );

    \I__5640\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26119\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__26122\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__26119\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5\
        );

    \I__5637\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26110\
        );

    \I__5636\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26107\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__26110\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__26107\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5\
        );

    \I__5633\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26099\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__26099\,
            I => \N__26096\
        );

    \I__5631\ : Span4Mux_v
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__5630\ : Odrv4
    port map (
            O => \N__26093\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_5\
        );

    \I__5629\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26084\
        );

    \I__5628\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26084\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__26084\,
            I => \N__26081\
        );

    \I__5626\ : Span4Mux_v
    port map (
            O => \N__26081\,
            I => \N__26078\
        );

    \I__5625\ : Odrv4
    port map (
            O => \N__26078\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_0\
        );

    \I__5624\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26071\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__26074\,
            I => \N__26068\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__26071\,
            I => \N__26065\
        );

    \I__5621\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26062\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__26065\,
            I => \N__26057\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26057\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__26057\,
            I => \N__26054\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__26054\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_4\
        );

    \I__5616\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26045\
        );

    \I__5615\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26045\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__5613\ : Span4Mux_v
    port map (
            O => \N__26042\,
            I => \N__26039\
        );

    \I__5612\ : Span4Mux_h
    port map (
            O => \N__26039\,
            I => \N__26036\
        );

    \I__5611\ : Odrv4
    port map (
            O => \N__26036\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_5\
        );

    \I__5610\ : InMux
    port map (
            O => \N__26033\,
            I => \N__26029\
        );

    \I__5609\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26026\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__26029\,
            I => \N__26023\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__26026\,
            I => \N__26020\
        );

    \I__5606\ : Span4Mux_h
    port map (
            O => \N__26023\,
            I => \N__26017\
        );

    \I__5605\ : Span4Mux_h
    port map (
            O => \N__26020\,
            I => \N__26014\
        );

    \I__5604\ : Odrv4
    port map (
            O => \N__26017\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1\
        );

    \I__5603\ : Odrv4
    port map (
            O => \N__26014\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1\
        );

    \I__5602\ : InMux
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__26006\,
            I => \N__26003\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__26003\,
            I => \N__25999\
        );

    \I__5599\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25996\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__25999\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__25996\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2\
        );

    \I__5596\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__25988\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_2\
        );

    \I__5594\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25982\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__25982\,
            I => \N__25978\
        );

    \I__5592\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25975\
        );

    \I__5591\ : Odrv4
    port map (
            O => \N__25978\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__25975\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3\
        );

    \I__5589\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__25967\,
            I => \N__25964\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__25964\,
            I => \N__25961\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__25961\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_3\
        );

    \I__5585\ : CEMux
    port map (
            O => \N__25958\,
            I => \N__25954\
        );

    \I__5584\ : CEMux
    port map (
            O => \N__25957\,
            I => \N__25951\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__25954\,
            I => \N__25948\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__25951\,
            I => \N__25945\
        );

    \I__5581\ : Span4Mux_v
    port map (
            O => \N__25948\,
            I => \N__25941\
        );

    \I__5580\ : Span4Mux_s3_v
    port map (
            O => \N__25945\,
            I => \N__25938\
        );

    \I__5579\ : CEMux
    port map (
            O => \N__25944\,
            I => \N__25935\
        );

    \I__5578\ : Span4Mux_h
    port map (
            O => \N__25941\,
            I => \N__25932\
        );

    \I__5577\ : Sp12to4
    port map (
            O => \N__25938\,
            I => \N__25929\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__25935\,
            I => \N__25926\
        );

    \I__5575\ : Sp12to4
    port map (
            O => \N__25932\,
            I => \N__25921\
        );

    \I__5574\ : Span12Mux_s8_h
    port map (
            O => \N__25929\,
            I => \N__25921\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__25926\,
            I => \N__25918\
        );

    \I__5572\ : Odrv12
    port map (
            O => \N__25921\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2\
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__25918\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2\
        );

    \I__5570\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25909\
        );

    \I__5569\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25906\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__25909\,
            I => \N__25903\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__25906\,
            I => \N__25900\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__25903\,
            I => \N__25897\
        );

    \I__5565\ : Span4Mux_h
    port map (
            O => \N__25900\,
            I => \N__25894\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__25897\,
            I => \N__25891\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__25894\,
            I => \N__25888\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__25891\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__25888\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0\
        );

    \I__5560\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25879\
        );

    \I__5559\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25876\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__25879\,
            I => \N__25873\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__25876\,
            I => \N__25870\
        );

    \I__5556\ : Span4Mux_h
    port map (
            O => \N__25873\,
            I => \N__25867\
        );

    \I__5555\ : Span4Mux_v
    port map (
            O => \N__25870\,
            I => \N__25864\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__25867\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1\
        );

    \I__5553\ : Odrv4
    port map (
            O => \N__25864\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1\
        );

    \I__5552\ : InMux
    port map (
            O => \N__25859\,
            I => \N__25856\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__25856\,
            I => \N__25853\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__25853\,
            I => \N__25850\
        );

    \I__5549\ : Span4Mux_s1_v
    port map (
            O => \N__25850\,
            I => \N__25846\
        );

    \I__5548\ : InMux
    port map (
            O => \N__25849\,
            I => \N__25843\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__25846\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__25843\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2\
        );

    \I__5545\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25835\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__5543\ : Odrv4
    port map (
            O => \N__25832\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_2\
        );

    \I__5542\ : CascadeMux
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__5541\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25823\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__25820\,
            I => \N__25817\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__25817\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_2\
        );

    \I__5537\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__25802\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_2\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__25799\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_2_cascade_\
        );

    \I__5531\ : SRMux
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__25793\,
            I => \N__25789\
        );

    \I__5529\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25786\
        );

    \I__5528\ : Span4Mux_h
    port map (
            O => \N__25789\,
            I => \N__25777\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__25786\,
            I => \N__25777\
        );

    \I__5526\ : InMux
    port map (
            O => \N__25785\,
            I => \N__25774\
        );

    \I__5525\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25770\
        );

    \I__5524\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25767\
        );

    \I__5523\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25764\
        );

    \I__5522\ : Span4Mux_v
    port map (
            O => \N__25777\,
            I => \N__25756\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__25774\,
            I => \N__25756\
        );

    \I__5520\ : InMux
    port map (
            O => \N__25773\,
            I => \N__25752\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__25770\,
            I => \N__25749\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__25767\,
            I => \N__25744\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__25764\,
            I => \N__25744\
        );

    \I__5516\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25741\
        );

    \I__5515\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25738\
        );

    \I__5514\ : InMux
    port map (
            O => \N__25761\,
            I => \N__25734\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__25756\,
            I => \N__25731\
        );

    \I__5512\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25728\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25725\
        );

    \I__5510\ : Span4Mux_v
    port map (
            O => \N__25749\,
            I => \N__25720\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__25744\,
            I => \N__25720\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__25741\,
            I => \N__25715\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__25738\,
            I => \N__25715\
        );

    \I__5506\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25712\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__25734\,
            I => \N__25709\
        );

    \I__5504\ : Span4Mux_v
    port map (
            O => \N__25731\,
            I => \N__25706\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__25728\,
            I => \N__25703\
        );

    \I__5502\ : Span4Mux_v
    port map (
            O => \N__25725\,
            I => \N__25700\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__25720\,
            I => \N__25693\
        );

    \I__5500\ : Span4Mux_v
    port map (
            O => \N__25715\,
            I => \N__25693\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__25712\,
            I => \N__25693\
        );

    \I__5498\ : Span12Mux_s9_h
    port map (
            O => \N__25709\,
            I => \N__25690\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__25706\,
            I => \N__25685\
        );

    \I__5496\ : Span4Mux_v
    port map (
            O => \N__25703\,
            I => \N__25685\
        );

    \I__5495\ : Span4Mux_s2_h
    port map (
            O => \N__25700\,
            I => \N__25680\
        );

    \I__5494\ : Span4Mux_h
    port map (
            O => \N__25693\,
            I => \N__25680\
        );

    \I__5493\ : Odrv12
    port map (
            O => \N__25690\,
            I => instruction_7
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__25685\,
            I => instruction_7
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__25680\,
            I => instruction_7
        );

    \I__5490\ : CascadeMux
    port map (
            O => \N__25673\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_2_cascade_\
        );

    \I__5489\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25662\
        );

    \I__5488\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25662\
        );

    \I__5487\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25653\
        );

    \I__5486\ : InMux
    port map (
            O => \N__25667\,
            I => \N__25653\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__25662\,
            I => \N__25650\
        );

    \I__5484\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25645\
        );

    \I__5483\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25645\
        );

    \I__5482\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25640\
        );

    \I__5481\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25640\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__25653\,
            I => \N__25632\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__25650\,
            I => \N__25627\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__25645\,
            I => \N__25627\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__25640\,
            I => \N__25624\
        );

    \I__5476\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25619\
        );

    \I__5475\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25619\
        );

    \I__5474\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25616\
        );

    \I__5473\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25613\
        );

    \I__5472\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25610\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__25632\,
            I => \N__25606\
        );

    \I__5470\ : Span4Mux_v
    port map (
            O => \N__25627\,
            I => \N__25598\
        );

    \I__5469\ : Span4Mux_v
    port map (
            O => \N__25624\,
            I => \N__25593\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__25619\,
            I => \N__25593\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__25616\,
            I => \N__25590\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__25613\,
            I => \N__25585\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__25610\,
            I => \N__25585\
        );

    \I__5464\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25582\
        );

    \I__5463\ : Span4Mux_v
    port map (
            O => \N__25606\,
            I => \N__25579\
        );

    \I__5462\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25574\
        );

    \I__5461\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25574\
        );

    \I__5460\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25571\
        );

    \I__5459\ : InMux
    port map (
            O => \N__25602\,
            I => \N__25566\
        );

    \I__5458\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25566\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__25598\,
            I => \N__25561\
        );

    \I__5456\ : Span4Mux_h
    port map (
            O => \N__25593\,
            I => \N__25561\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__25590\,
            I => \N__25556\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__25585\,
            I => \N__25556\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__25582\,
            I => \processor_zipi8.bank\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__25579\,
            I => \processor_zipi8.bank\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__25574\,
            I => \processor_zipi8.bank\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__25571\,
            I => \processor_zipi8.bank\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__25566\,
            I => \processor_zipi8.bank\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__25561\,
            I => \processor_zipi8.bank\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__25556\,
            I => \processor_zipi8.bank\
        );

    \I__5446\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25537\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__25540\,
            I => \N__25534\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__25537\,
            I => \N__25531\
        );

    \I__5443\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25528\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__25531\,
            I => \N__25525\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__25528\,
            I => \N__25522\
        );

    \I__5440\ : Span4Mux_v
    port map (
            O => \N__25525\,
            I => \N__25517\
        );

    \I__5439\ : Span4Mux_s3_h
    port map (
            O => \N__25522\,
            I => \N__25517\
        );

    \I__5438\ : Span4Mux_s3_v
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__25514\,
            I => \N__25511\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__25511\,
            I => \processor_zipi8.sy_2\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__25508\,
            I => \N__25505\
        );

    \I__5434\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25501\
        );

    \I__5433\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25498\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__25501\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__25498\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2\
        );

    \I__5430\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25490\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__25490\,
            I => \N__25486\
        );

    \I__5428\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__25486\,
            I => \N__25480\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__25483\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__25480\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__25475\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_2_cascade_\
        );

    \I__5423\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25469\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__25469\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_2\
        );

    \I__5421\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25460\
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__25460\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_2\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__25457\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_2_cascade_\
        );

    \I__5417\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25451\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__25451\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_2\
        );

    \I__5415\ : InMux
    port map (
            O => \N__25448\,
            I => \N__25444\
        );

    \I__5414\ : InMux
    port map (
            O => \N__25447\,
            I => \N__25441\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__25444\,
            I => \N__25438\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__25441\,
            I => \N__25435\
        );

    \I__5411\ : Span4Mux_v
    port map (
            O => \N__25438\,
            I => \N__25430\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__25435\,
            I => \N__25430\
        );

    \I__5409\ : Span4Mux_v
    port map (
            O => \N__25430\,
            I => \N__25427\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__25427\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_0\
        );

    \I__5407\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25420\
        );

    \I__5406\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25417\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__25420\,
            I => \N__25414\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__25417\,
            I => \N__25411\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__25414\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1\
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__25411\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__25406\,
            I => \N__25402\
        );

    \I__5400\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25399\
        );

    \I__5399\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25396\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__25399\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__25396\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1\
        );

    \I__5396\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25387\
        );

    \I__5395\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25384\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__25387\,
            I => \N__25379\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__25384\,
            I => \N__25379\
        );

    \I__5392\ : Span4Mux_h
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__25376\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_1\
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__25373\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_1_cascade_\
        );

    \I__5389\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25366\
        );

    \I__5388\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25363\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__25366\,
            I => \N__25358\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__25363\,
            I => \N__25358\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__25355\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_1\
        );

    \I__5383\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25349\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__25349\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1\
        );

    \I__5381\ : CEMux
    port map (
            O => \N__25346\,
            I => \N__25343\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__25343\,
            I => \N__25340\
        );

    \I__5379\ : Span4Mux_h
    port map (
            O => \N__25340\,
            I => \N__25336\
        );

    \I__5378\ : CEMux
    port map (
            O => \N__25339\,
            I => \N__25331\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__25336\,
            I => \N__25328\
        );

    \I__5376\ : CEMux
    port map (
            O => \N__25335\,
            I => \N__25325\
        );

    \I__5375\ : CEMux
    port map (
            O => \N__25334\,
            I => \N__25322\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__25331\,
            I => \N__25319\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__25328\,
            I => \N__25314\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__25325\,
            I => \N__25314\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25311\
        );

    \I__5370\ : Span4Mux_v
    port map (
            O => \N__25319\,
            I => \N__25308\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__25314\,
            I => \N__25305\
        );

    \I__5368\ : Sp12to4
    port map (
            O => \N__25311\,
            I => \N__25302\
        );

    \I__5367\ : Span4Mux_s0_h
    port map (
            O => \N__25308\,
            I => \N__25299\
        );

    \I__5366\ : IoSpan4Mux
    port map (
            O => \N__25305\,
            I => \N__25296\
        );

    \I__5365\ : Span12Mux_v
    port map (
            O => \N__25302\,
            I => \N__25291\
        );

    \I__5364\ : Sp12to4
    port map (
            O => \N__25299\,
            I => \N__25291\
        );

    \I__5363\ : Span4Mux_s3_v
    port map (
            O => \N__25296\,
            I => \N__25288\
        );

    \I__5362\ : Odrv12
    port map (
            O => \N__25291\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__25288\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0\
        );

    \I__5360\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25279\
        );

    \I__5359\ : InMux
    port map (
            O => \N__25282\,
            I => \N__25276\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__25279\,
            I => \N__25273\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__25276\,
            I => \N__25270\
        );

    \I__5356\ : Span4Mux_h
    port map (
            O => \N__25273\,
            I => \N__25265\
        );

    \I__5355\ : Span4Mux_s3_h
    port map (
            O => \N__25270\,
            I => \N__25265\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__25265\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_4\
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__25262\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_4_cascade_\
        );

    \I__5352\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25256\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__25253\,
            I => \N__25249\
        );

    \I__5349\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25246\
        );

    \I__5348\ : Odrv4
    port map (
            O => \N__25249\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__25246\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__25241\,
            I => \N__25238\
        );

    \I__5345\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25234\
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__25237\,
            I => \N__25231\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__25234\,
            I => \N__25228\
        );

    \I__5342\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25225\
        );

    \I__5341\ : Odrv12
    port map (
            O => \N__25228\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__25225\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4\
        );

    \I__5339\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25217\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__25217\,
            I => \N__25213\
        );

    \I__5337\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25210\
        );

    \I__5336\ : Span4Mux_v
    port map (
            O => \N__25213\,
            I => \N__25205\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__25210\,
            I => \N__25205\
        );

    \I__5334\ : Span4Mux_v
    port map (
            O => \N__25205\,
            I => \N__25202\
        );

    \I__5333\ : Span4Mux_s1_v
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__25199\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_4\
        );

    \I__5331\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25192\
        );

    \I__5330\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25189\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__25192\,
            I => \N__25186\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__25189\,
            I => \N__25183\
        );

    \I__5327\ : Span12Mux_v
    port map (
            O => \N__25186\,
            I => \N__25180\
        );

    \I__5326\ : Span4Mux_h
    port map (
            O => \N__25183\,
            I => \N__25177\
        );

    \I__5325\ : Odrv12
    port map (
            O => \N__25180\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__25177\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__25172\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_4_cascade_\
        );

    \I__5322\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__25166\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_4\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__25163\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_4_cascade_\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__25160\,
            I => \N__25157\
        );

    \I__5318\ : InMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__25154\,
            I => \N__25151\
        );

    \I__5316\ : Odrv12
    port map (
            O => \N__25151\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_4\
        );

    \I__5315\ : CascadeMux
    port map (
            O => \N__25148\,
            I => \N__25144\
        );

    \I__5314\ : InMux
    port map (
            O => \N__25147\,
            I => \N__25139\
        );

    \I__5313\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25139\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__25139\,
            I => \N__25136\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__25136\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_4\
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__25133\,
            I => \N__25130\
        );

    \I__5309\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25124\
        );

    \I__5308\ : InMux
    port map (
            O => \N__25129\,
            I => \N__25124\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__25124\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_4\
        );

    \I__5306\ : CascadeMux
    port map (
            O => \N__25121\,
            I => \N__25118\
        );

    \I__5305\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__5303\ : Odrv4
    port map (
            O => \N__25112\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_4\
        );

    \I__5302\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25105\
        );

    \I__5301\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25102\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__25105\,
            I => \N__25097\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__25102\,
            I => \N__25097\
        );

    \I__5298\ : Span4Mux_h
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__5297\ : Odrv4
    port map (
            O => \N__25094\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_4\
        );

    \I__5296\ : CEMux
    port map (
            O => \N__25091\,
            I => \N__25088\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__25088\,
            I => \N__25084\
        );

    \I__5294\ : CEMux
    port map (
            O => \N__25087\,
            I => \N__25081\
        );

    \I__5293\ : Span4Mux_v
    port map (
            O => \N__25084\,
            I => \N__25078\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25075\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__25078\,
            I => \N__25072\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__25075\,
            I => \N__25069\
        );

    \I__5289\ : Sp12to4
    port map (
            O => \N__25072\,
            I => \N__25064\
        );

    \I__5288\ : Sp12to4
    port map (
            O => \N__25069\,
            I => \N__25064\
        );

    \I__5287\ : Odrv12
    port map (
            O => \N__25064\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe16\
        );

    \I__5286\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25058\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__25058\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__5283\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__25049\,
            I => \N__25045\
        );

    \I__5281\ : InMux
    port map (
            O => \N__25048\,
            I => \N__25042\
        );

    \I__5280\ : Span4Mux_h
    port map (
            O => \N__25045\,
            I => \N__25039\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__25042\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__25039\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5\
        );

    \I__5277\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25030\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__25033\,
            I => \N__25027\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__25024\
        );

    \I__5274\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25021\
        );

    \I__5273\ : Span4Mux_v
    port map (
            O => \N__25024\,
            I => \N__25018\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__25021\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__25018\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5\
        );

    \I__5270\ : CascadeMux
    port map (
            O => \N__25013\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_5_cascade_\
        );

    \I__5269\ : InMux
    port map (
            O => \N__25010\,
            I => \N__25007\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__5267\ : Span4Mux_s3_h
    port map (
            O => \N__25004\,
            I => \N__25001\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__25001\,
            I => \N__24998\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__24998\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_5\
        );

    \I__5264\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__24992\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_5\
        );

    \I__5262\ : CascadeMux
    port map (
            O => \N__24989\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_5_cascade_\
        );

    \I__5261\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__24980\,
            I => \N__24977\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__24974\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_5\
        );

    \I__5256\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24968\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__24968\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_1\
        );

    \I__5254\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24962\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__24962\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_1\
        );

    \I__5252\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__24956\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_1\
        );

    \I__5250\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24947\
        );

    \I__5249\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24947\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__24947\,
            I => \N__24944\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__24944\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_4\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__24941\,
            I => \N__24937\
        );

    \I__5245\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24934\
        );

    \I__5244\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24931\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__24934\,
            I => \N__24928\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__24931\,
            I => \N__24925\
        );

    \I__5241\ : Span4Mux_v
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__24925\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__24922\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5\
        );

    \I__5238\ : CEMux
    port map (
            O => \N__24917\,
            I => \N__24913\
        );

    \I__5237\ : CEMux
    port map (
            O => \N__24916\,
            I => \N__24910\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__24913\,
            I => \N__24907\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__24910\,
            I => \N__24904\
        );

    \I__5234\ : Span4Mux_s2_v
    port map (
            O => \N__24907\,
            I => \N__24901\
        );

    \I__5233\ : Span12Mux_s8_h
    port map (
            O => \N__24904\,
            I => \N__24898\
        );

    \I__5232\ : Span4Mux_h
    port map (
            O => \N__24901\,
            I => \N__24895\
        );

    \I__5231\ : Odrv12
    port map (
            O => \N__24898\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__24895\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17\
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__24890\,
            I => \N__24887\
        );

    \I__5228\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24884\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__24884\,
            I => \N__24881\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__24881\,
            I => \N__24878\
        );

    \I__5225\ : Span4Mux_s3_h
    port map (
            O => \N__24878\,
            I => \N__24874\
        );

    \I__5224\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24871\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__24874\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__24871\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6\
        );

    \I__5221\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24859\
        );

    \I__5219\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24856\
        );

    \I__5218\ : Span4Mux_v
    port map (
            O => \N__24859\,
            I => \N__24851\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__24856\,
            I => \N__24851\
        );

    \I__5216\ : Span4Mux_v
    port map (
            O => \N__24851\,
            I => \N__24848\
        );

    \I__5215\ : Odrv4
    port map (
            O => \N__24848\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_6\
        );

    \I__5214\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__5212\ : Odrv12
    port map (
            O => \N__24839\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_6\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__5210\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24829\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__24832\,
            I => \N__24826\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24823\
        );

    \I__5207\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24820\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__24823\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__24820\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0\
        );

    \I__5204\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__5203\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24805\
        );

    \I__5201\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24802\
        );

    \I__5200\ : Span4Mux_v
    port map (
            O => \N__24805\,
            I => \N__24799\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__24802\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__24799\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__24794\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_0_cascade_\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__24791\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI86UU1_0_cascade_\
        );

    \I__5195\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__24785\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNI2KHQ1_0\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__24782\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_0_cascade_\
        );

    \I__5192\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24776\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__5190\ : Span4Mux_v
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__5189\ : Span4Mux_h
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__24767\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFG9I8_0\
        );

    \I__5187\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24761\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24757\
        );

    \I__5185\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24754\
        );

    \I__5184\ : Span4Mux_s3_h
    port map (
            O => \N__24757\,
            I => \N__24751\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__24754\,
            I => \N__24748\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__24751\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0\
        );

    \I__5181\ : Odrv12
    port map (
            O => \N__24748\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__24743\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_0_cascade_\
        );

    \I__5179\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24737\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__24737\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIKPJ32_0\
        );

    \I__5177\ : InMux
    port map (
            O => \N__24734\,
            I => \N__24731\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__5175\ : Odrv4
    port map (
            O => \N__24728\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_0\
        );

    \I__5174\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24722\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__24722\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI4QLM1_0\
        );

    \I__5172\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24715\
        );

    \I__5171\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24712\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__24715\,
            I => \N__24709\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__24712\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0\
        );

    \I__5168\ : Odrv12
    port map (
            O => \N__24709\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0\
        );

    \I__5167\ : CascadeMux
    port map (
            O => \N__24704\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_0_cascade_\
        );

    \I__5166\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24698\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__24695\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_0\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__24692\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_0_cascade_\
        );

    \I__5162\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24686\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__24686\,
            I => \N__24683\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__24683\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_0\
        );

    \I__5159\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24677\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__24677\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_0\
        );

    \I__5157\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__24671\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_0\
        );

    \I__5155\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24662\
        );

    \I__5154\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24662\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__24662\,
            I => \N__24659\
        );

    \I__5152\ : Odrv12
    port map (
            O => \N__24659\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_0\
        );

    \I__5151\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24653\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__24653\,
            I => \N__24649\
        );

    \I__5149\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24646\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__24649\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__24646\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0\
        );

    \I__5146\ : CascadeMux
    port map (
            O => \N__24641\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_0_cascade_\
        );

    \I__5145\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__24632\,
            I => \N__24628\
        );

    \I__5142\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24625\
        );

    \I__5141\ : Odrv4
    port map (
            O => \N__24628\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__24625\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0\
        );

    \I__5139\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__24614\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_6\
        );

    \I__5136\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__24605\,
            I => \N__24602\
        );

    \I__5133\ : Span4Mux_h
    port map (
            O => \N__24602\,
            I => \N__24599\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__24599\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_6\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__24596\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_4_cascade_\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__24593\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_4_cascade_\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__24590\,
            I => \N__24587\
        );

    \I__5128\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__24581\,
            I => \N__24578\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__24578\,
            I => \N__24575\
        );

    \I__5124\ : Odrv4
    port map (
            O => \N__24575\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_4\
        );

    \I__5123\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24568\
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__24571\,
            I => \N__24565\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24562\
        );

    \I__5120\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24559\
        );

    \I__5119\ : Span4Mux_s3_v
    port map (
            O => \N__24562\,
            I => \N__24554\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__24559\,
            I => \N__24554\
        );

    \I__5117\ : Span4Mux_v
    port map (
            O => \N__24554\,
            I => \N__24551\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__24551\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_6\
        );

    \I__5115\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24544\
        );

    \I__5114\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24541\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__24544\,
            I => \N__24538\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__24541\,
            I => \N__24535\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__24538\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6\
        );

    \I__5110\ : Odrv12
    port map (
            O => \N__24535\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__5108\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__24524\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_6\
        );

    \I__5106\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24514\
        );

    \I__5104\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24511\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__24514\,
            I => \N__24508\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__24511\,
            I => \N__24505\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__24508\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__24505\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4\
        );

    \I__5099\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24496\
        );

    \I__5098\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24493\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__24496\,
            I => \N__24490\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__24493\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__24490\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4\
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__24485\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_4_cascade_\
        );

    \I__5093\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24475\
        );

    \I__5091\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24472\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__24475\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__24472\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4\
        );

    \I__5088\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__24464\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_4\
        );

    \I__5086\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24458\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__24458\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_6\
        );

    \I__5084\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24452\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__24452\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_6\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__5081\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24440\
        );

    \I__5080\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24440\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__24440\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_6\
        );

    \I__5078\ : CEMux
    port map (
            O => \N__24437\,
            I => \N__24434\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__24431\,
            I => \N__24428\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__24428\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe28\
        );

    \I__5074\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24421\
        );

    \I__5073\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24418\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__24421\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__24418\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5\
        );

    \I__5070\ : CEMux
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__24410\,
            I => \N__24405\
        );

    \I__5068\ : CEMux
    port map (
            O => \N__24409\,
            I => \N__24402\
        );

    \I__5067\ : CEMux
    port map (
            O => \N__24408\,
            I => \N__24399\
        );

    \I__5066\ : Span4Mux_s3_v
    port map (
            O => \N__24405\,
            I => \N__24394\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__24402\,
            I => \N__24394\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__24399\,
            I => \N__24391\
        );

    \I__5063\ : Span4Mux_v
    port map (
            O => \N__24394\,
            I => \N__24388\
        );

    \I__5062\ : Span4Mux_v
    port map (
            O => \N__24391\,
            I => \N__24385\
        );

    \I__5061\ : Span4Mux_h
    port map (
            O => \N__24388\,
            I => \N__24382\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__24385\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__24382\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30\
        );

    \I__5058\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24374\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__24374\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_6\
        );

    \I__5056\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24368\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__24368\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_6\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__24365\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_6_cascade_\
        );

    \I__5053\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24356\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__24356\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNISIMM1_6\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__24353\,
            I => \N__24349\
        );

    \I__5049\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24344\
        );

    \I__5048\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24344\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__24344\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_5\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__24341\,
            I => \N__24334\
        );

    \I__5045\ : CascadeMux
    port map (
            O => \N__24340\,
            I => \N__24328\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__24339\,
            I => \N__24324\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__24338\,
            I => \N__24320\
        );

    \I__5042\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24311\
        );

    \I__5041\ : InMux
    port map (
            O => \N__24334\,
            I => \N__24301\
        );

    \I__5040\ : InMux
    port map (
            O => \N__24333\,
            I => \N__24301\
        );

    \I__5039\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24301\
        );

    \I__5038\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24294\
        );

    \I__5037\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24294\
        );

    \I__5036\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24294\
        );

    \I__5035\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24279\
        );

    \I__5034\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24279\
        );

    \I__5033\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24279\
        );

    \I__5032\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24279\
        );

    \I__5031\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24272\
        );

    \I__5030\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24267\
        );

    \I__5029\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24267\
        );

    \I__5028\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24264\
        );

    \I__5027\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24261\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__24311\,
            I => \N__24258\
        );

    \I__5025\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24255\
        );

    \I__5024\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24250\
        );

    \I__5023\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24250\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__24301\,
            I => \N__24245\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24245\
        );

    \I__5020\ : InMux
    port map (
            O => \N__24293\,
            I => \N__24240\
        );

    \I__5019\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24240\
        );

    \I__5018\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24237\
        );

    \I__5017\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24230\
        );

    \I__5016\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24230\
        );

    \I__5015\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24230\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__24279\,
            I => \N__24227\
        );

    \I__5013\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24218\
        );

    \I__5012\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24218\
        );

    \I__5011\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24218\
        );

    \I__5010\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24218\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__24272\,
            I => \N__24215\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__24267\,
            I => \N__24212\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__24264\,
            I => \N__24203\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__24261\,
            I => \N__24203\
        );

    \I__5005\ : Span4Mux_h
    port map (
            O => \N__24258\,
            I => \N__24203\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__24255\,
            I => \N__24203\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__24250\,
            I => \N__24194\
        );

    \I__5002\ : Span4Mux_h
    port map (
            O => \N__24245\,
            I => \N__24194\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24194\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__24237\,
            I => \N__24194\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24187\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__24227\,
            I => \N__24187\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24187\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__24215\,
            I => \N__24178\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__24212\,
            I => \N__24178\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__24203\,
            I => \N__24178\
        );

    \I__4993\ : Span4Mux_v
    port map (
            O => \N__24194\,
            I => \N__24178\
        );

    \I__4992\ : Odrv4
    port map (
            O => \N__24187\,
            I => instruction_16
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__24178\,
            I => instruction_16
        );

    \I__4990\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24156\
        );

    \I__4989\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24156\
        );

    \I__4988\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24148\
        );

    \I__4987\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24148\
        );

    \I__4986\ : CascadeMux
    port map (
            O => \N__24169\,
            I => \N__24144\
        );

    \I__4985\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24139\
        );

    \I__4984\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24139\
        );

    \I__4983\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24136\
        );

    \I__4982\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24127\
        );

    \I__4981\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24127\
        );

    \I__4980\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24127\
        );

    \I__4979\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24127\
        );

    \I__4978\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24123\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__24156\,
            I => \N__24120\
        );

    \I__4976\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24113\
        );

    \I__4975\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24113\
        );

    \I__4974\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24113\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__24148\,
            I => \N__24108\
        );

    \I__4972\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24105\
        );

    \I__4971\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24102\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__24139\,
            I => \N__24091\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__24136\,
            I => \N__24086\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24086\
        );

    \I__4967\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24083\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__24123\,
            I => \N__24076\
        );

    \I__4965\ : Span4Mux_s3_v
    port map (
            O => \N__24120\,
            I => \N__24076\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__24113\,
            I => \N__24076\
        );

    \I__4963\ : InMux
    port map (
            O => \N__24112\,
            I => \N__24073\
        );

    \I__4962\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24070\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__24108\,
            I => \N__24063\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24063\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24063\
        );

    \I__4958\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24054\
        );

    \I__4957\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24054\
        );

    \I__4956\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24054\
        );

    \I__4955\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24054\
        );

    \I__4954\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24045\
        );

    \I__4953\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24045\
        );

    \I__4952\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24045\
        );

    \I__4951\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24045\
        );

    \I__4950\ : Span4Mux_s3_v
    port map (
            O => \N__24091\,
            I => \N__24036\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__24086\,
            I => \N__24036\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__24083\,
            I => \N__24036\
        );

    \I__4947\ : Span4Mux_h
    port map (
            O => \N__24076\,
            I => \N__24036\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__24073\,
            I => \N__24025\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__24025\
        );

    \I__4944\ : Sp12to4
    port map (
            O => \N__24063\,
            I => \N__24025\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24025\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__24025\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__24036\,
            I => \N__24022\
        );

    \I__4940\ : Span12Mux_s9_h
    port map (
            O => \N__24025\,
            I => \N__24019\
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__24022\,
            I => instruction_15
        );

    \I__4938\ : Odrv12
    port map (
            O => \N__24019\,
            I => instruction_15
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__24014\,
            I => \N__24009\
        );

    \I__4936\ : InMux
    port map (
            O => \N__24013\,
            I => \N__24006\
        );

    \I__4935\ : InMux
    port map (
            O => \N__24012\,
            I => \N__24003\
        );

    \I__4934\ : InMux
    port map (
            O => \N__24009\,
            I => \N__24000\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__24006\,
            I => \N__23994\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__24003\,
            I => \N__23994\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__24000\,
            I => \N__23991\
        );

    \I__4930\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23982\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__23994\,
            I => \N__23977\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__23991\,
            I => \N__23977\
        );

    \I__4927\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23971\
        );

    \I__4926\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23971\
        );

    \I__4925\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23968\
        );

    \I__4924\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23965\
        );

    \I__4923\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23962\
        );

    \I__4922\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23959\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__23982\,
            I => \N__23956\
        );

    \I__4920\ : IoSpan4Mux
    port map (
            O => \N__23977\,
            I => \N__23953\
        );

    \I__4919\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23950\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__23971\,
            I => \N__23947\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__23968\,
            I => \N__23944\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__23965\,
            I => \N__23941\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__23962\,
            I => \N__23938\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23935\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__23956\,
            I => \N__23932\
        );

    \I__4912\ : Span4Mux_s3_h
    port map (
            O => \N__23953\,
            I => \N__23927\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__23950\,
            I => \N__23927\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__23947\,
            I => \N__23922\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__23944\,
            I => \N__23922\
        );

    \I__4908\ : Span4Mux_h
    port map (
            O => \N__23941\,
            I => \N__23919\
        );

    \I__4907\ : Span12Mux_s7_h
    port map (
            O => \N__23938\,
            I => \N__23916\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__23935\,
            I => \N__23913\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__23932\,
            I => \N__23908\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__23927\,
            I => \N__23908\
        );

    \I__4903\ : Span4Mux_v
    port map (
            O => \N__23922\,
            I => \N__23905\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__23919\,
            I => \processor_zipi8.un28_carry_flag_value_1\
        );

    \I__4901\ : Odrv12
    port map (
            O => \N__23916\,
            I => \processor_zipi8.un28_carry_flag_value_1\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__23913\,
            I => \processor_zipi8.un28_carry_flag_value_1\
        );

    \I__4899\ : Odrv4
    port map (
            O => \N__23908\,
            I => \processor_zipi8.un28_carry_flag_value_1\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__23905\,
            I => \processor_zipi8.un28_carry_flag_value_1\
        );

    \I__4897\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__23891\,
            I => \N__23887\
        );

    \I__4895\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23884\
        );

    \I__4894\ : Span4Mux_h
    port map (
            O => \N__23887\,
            I => \N__23879\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__23884\,
            I => \N__23879\
        );

    \I__4892\ : Span4Mux_v
    port map (
            O => \N__23879\,
            I => \N__23876\
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__23876\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_5\
        );

    \I__4890\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23869\
        );

    \I__4889\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23866\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__23869\,
            I => \N__23863\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__23866\,
            I => \N__23860\
        );

    \I__4886\ : Span4Mux_h
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__23860\,
            I => \N__23854\
        );

    \I__4884\ : Span4Mux_v
    port map (
            O => \N__23857\,
            I => \N__23851\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__23854\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__23851\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7\
        );

    \I__4881\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__23843\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_6\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__23840\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_6_cascade_\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23834\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__23834\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_6\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__23831\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_6_cascade_\
        );

    \I__4875\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23825\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__23825\,
            I => \N__23822\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__23822\,
            I => \N__23819\
        );

    \I__4872\ : Span4Mux_h
    port map (
            O => \N__23819\,
            I => \N__23816\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__23816\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_6\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__4869\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23806\
        );

    \I__4868\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23803\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__23806\,
            I => \N__23798\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__23803\,
            I => \N__23798\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__23798\,
            I => \N__23795\
        );

    \I__4864\ : Span4Mux_v
    port map (
            O => \N__23795\,
            I => \N__23792\
        );

    \I__4863\ : Span4Mux_v
    port map (
            O => \N__23792\,
            I => \N__23789\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__23789\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_6\
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__23786\,
            I => \N__23783\
        );

    \I__4860\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23777\
        );

    \I__4859\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23777\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__23777\,
            I => \N__23774\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__23774\,
            I => \N__23771\
        );

    \I__4856\ : Sp12to4
    port map (
            O => \N__23771\,
            I => \N__23768\
        );

    \I__4855\ : Span12Mux_v
    port map (
            O => \N__23768\,
            I => \N__23765\
        );

    \I__4854\ : Odrv12
    port map (
            O => \N__23765\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_7\
        );

    \I__4853\ : CEMux
    port map (
            O => \N__23762\,
            I => \N__23759\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__23759\,
            I => \N__23756\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__4850\ : Span4Mux_v
    port map (
            O => \N__23753\,
            I => \N__23750\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__23750\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe1\
        );

    \I__4848\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__23744\,
            I => \N__23740\
        );

    \I__4846\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23737\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__23740\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__23737\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__23732\,
            I => \N__23729\
        );

    \I__4842\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23726\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__23726\,
            I => \N__23723\
        );

    \I__4840\ : Span4Mux_s2_v
    port map (
            O => \N__23723\,
            I => \N__23719\
        );

    \I__4839\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23716\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__23719\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__23716\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5\
        );

    \I__4836\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__4834\ : Span4Mux_h
    port map (
            O => \N__23705\,
            I => \N__23701\
        );

    \I__4833\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23698\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__23701\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__23698\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__23693\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_5_cascade_\
        );

    \I__4829\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__23687\,
            I => \N__23683\
        );

    \I__4827\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23680\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__23683\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__23680\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__23675\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_5_cascade_\
        );

    \I__4823\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__23669\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_123\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__23666\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_99_cascade_\
        );

    \I__4820\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__4818\ : Span4Mux_s3_h
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__4817\ : Span4Mux_h
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__23651\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_5\
        );

    \I__4815\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__4812\ : Span4Mux_h
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__23636\,
            I => \processor_zipi8.stack_memory_3\
        );

    \I__4810\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__4808\ : Span4Mux_h
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__23624\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_3\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__4805\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__4803\ : Span4Mux_v
    port map (
            O => \N__23612\,
            I => \N__23608\
        );

    \I__4802\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23605\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__23608\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__23605\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3\
        );

    \I__4799\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23597\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__23597\,
            I => \N__23593\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__23596\,
            I => \N__23590\
        );

    \I__4796\ : Span4Mux_s3_v
    port map (
            O => \N__23593\,
            I => \N__23587\
        );

    \I__4795\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23584\
        );

    \I__4794\ : Odrv4
    port map (
            O => \N__23587\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__23584\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3\
        );

    \I__4792\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__4790\ : Odrv4
    port map (
            O => \N__23573\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_3\
        );

    \I__4789\ : CEMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__4787\ : Span4Mux_h
    port map (
            O => \N__23564\,
            I => \N__23560\
        );

    \I__4786\ : CEMux
    port map (
            O => \N__23563\,
            I => \N__23557\
        );

    \I__4785\ : Span4Mux_s1_h
    port map (
            O => \N__23560\,
            I => \N__23554\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__23557\,
            I => \N__23551\
        );

    \I__4783\ : Sp12to4
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__23551\,
            I => \N__23545\
        );

    \I__4781\ : Span12Mux_v
    port map (
            O => \N__23548\,
            I => \N__23542\
        );

    \I__4780\ : Sp12to4
    port map (
            O => \N__23545\,
            I => \N__23539\
        );

    \I__4779\ : Odrv12
    port map (
            O => \N__23542\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4\
        );

    \I__4778\ : Odrv12
    port map (
            O => \N__23539\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4\
        );

    \I__4777\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23530\
        );

    \I__4776\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23527\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__23530\,
            I => \N__23524\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__4773\ : Span4Mux_v
    port map (
            O => \N__23524\,
            I => \N__23518\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__23521\,
            I => \N__23515\
        );

    \I__4771\ : Odrv4
    port map (
            O => \N__23518\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__23515\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0\
        );

    \I__4769\ : CascadeMux
    port map (
            O => \N__23510\,
            I => \N__23506\
        );

    \I__4768\ : CascadeMux
    port map (
            O => \N__23509\,
            I => \N__23503\
        );

    \I__4767\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23500\
        );

    \I__4766\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23497\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__23500\,
            I => \N__23494\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__23497\,
            I => \N__23491\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__23494\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1\
        );

    \I__4762\ : Odrv12
    port map (
            O => \N__23491\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__23486\,
            I => \N__23482\
        );

    \I__4760\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23479\
        );

    \I__4759\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23476\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23473\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__23476\,
            I => \N__23470\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__23473\,
            I => \N__23467\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__23470\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3\
        );

    \I__4754\ : Odrv4
    port map (
            O => \N__23467\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3\
        );

    \I__4753\ : CascadeMux
    port map (
            O => \N__23462\,
            I => \N__23458\
        );

    \I__4752\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23455\
        );

    \I__4751\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23452\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__23455\,
            I => \N__23447\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__23452\,
            I => \N__23447\
        );

    \I__4748\ : Sp12to4
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__4747\ : Span12Mux_s11_v
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__4746\ : Odrv12
    port map (
            O => \N__23441\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_6\
        );

    \I__4745\ : CEMux
    port map (
            O => \N__23438\,
            I => \N__23434\
        );

    \I__4744\ : CEMux
    port map (
            O => \N__23437\,
            I => \N__23431\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__23434\,
            I => \N__23428\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N__23425\
        );

    \I__4741\ : Span4Mux_v
    port map (
            O => \N__23428\,
            I => \N__23422\
        );

    \I__4740\ : Span4Mux_s0_v
    port map (
            O => \N__23425\,
            I => \N__23419\
        );

    \I__4739\ : Span4Mux_v
    port map (
            O => \N__23422\,
            I => \N__23416\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__23419\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5\
        );

    \I__4737\ : Odrv4
    port map (
            O => \N__23416\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5\
        );

    \I__4736\ : InMux
    port map (
            O => \N__23411\,
            I => \N__23408\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__23408\,
            I => \N__23404\
        );

    \I__4734\ : InMux
    port map (
            O => \N__23407\,
            I => \N__23401\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__23404\,
            I => \N__23398\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__23401\,
            I => \N__23395\
        );

    \I__4731\ : Span4Mux_v
    port map (
            O => \N__23398\,
            I => \N__23390\
        );

    \I__4730\ : Span4Mux_h
    port map (
            O => \N__23395\,
            I => \N__23390\
        );

    \I__4729\ : Odrv4
    port map (
            O => \N__23390\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_0\
        );

    \I__4728\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23383\
        );

    \I__4727\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23380\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__23383\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__23380\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2\
        );

    \I__4724\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23372\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__23372\,
            I => \N__23368\
        );

    \I__4722\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23365\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__23368\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__23365\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2\
        );

    \I__4719\ : CascadeMux
    port map (
            O => \N__23360\,
            I => \N__23356\
        );

    \I__4718\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23351\
        );

    \I__4717\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23351\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__4714\ : Sp12to4
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__4713\ : Odrv12
    port map (
            O => \N__23342\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_4\
        );

    \I__4712\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23335\
        );

    \I__4711\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23332\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__23335\,
            I => \N__23329\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__23332\,
            I => \N__23326\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__23329\,
            I => \N__23323\
        );

    \I__4707\ : Span12Mux_s10_v
    port map (
            O => \N__23326\,
            I => \N__23320\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__23323\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5\
        );

    \I__4705\ : Odrv12
    port map (
            O => \N__23320\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5\
        );

    \I__4704\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23308\
        );

    \I__4702\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23305\
        );

    \I__4701\ : Span4Mux_v
    port map (
            O => \N__23308\,
            I => \N__23302\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__23305\,
            I => \N__23299\
        );

    \I__4699\ : Span4Mux_v
    port map (
            O => \N__23302\,
            I => \N__23294\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__23299\,
            I => \N__23294\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__23294\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_7\
        );

    \I__4696\ : CEMux
    port map (
            O => \N__23291\,
            I => \N__23288\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__23288\,
            I => \N__23285\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__23285\,
            I => \N__23282\
        );

    \I__4693\ : Span4Mux_h
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__4692\ : Odrv4
    port map (
            O => \N__23279\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe23\
        );

    \I__4691\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23272\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__23275\,
            I => \N__23269\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__23272\,
            I => \N__23266\
        );

    \I__4688\ : InMux
    port map (
            O => \N__23269\,
            I => \N__23263\
        );

    \I__4687\ : Span4Mux_v
    port map (
            O => \N__23266\,
            I => \N__23258\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__23263\,
            I => \N__23258\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__23258\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_0\
        );

    \I__4684\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23252\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__23252\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_1_0\
        );

    \I__4682\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23245\
        );

    \I__4681\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23242\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23237\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__23242\,
            I => \N__23237\
        );

    \I__4678\ : Span4Mux_v
    port map (
            O => \N__23237\,
            I => \N__23234\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__23234\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_1\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__23231\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_1_cascade_\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__23228\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_cascade_\
        );

    \I__4674\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__23219\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__23216\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_cascade_\
        );

    \I__4670\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__23210\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__23207\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_cascade_\
        );

    \I__4667\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23201\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__23201\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_1\
        );

    \I__4665\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__23195\,
            I => \N__23192\
        );

    \I__4663\ : Span4Mux_v
    port map (
            O => \N__23192\,
            I => \N__23188\
        );

    \I__4662\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23185\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__23188\,
            I => \processor_zipi8.sy_1\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__23185\,
            I => \processor_zipi8.sy_1\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__23180\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_4_cascade_\
        );

    \I__4658\ : InMux
    port map (
            O => \N__23177\,
            I => \N__23174\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__4656\ : Span4Mux_v
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__23168\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNICSGN1_4\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__23165\,
            I => \N__23160\
        );

    \I__4653\ : CascadeMux
    port map (
            O => \N__23164\,
            I => \N__23155\
        );

    \I__4652\ : CascadeMux
    port map (
            O => \N__23163\,
            I => \N__23150\
        );

    \I__4651\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23147\
        );

    \I__4650\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23133\
        );

    \I__4649\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23133\
        );

    \I__4648\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23133\
        );

    \I__4647\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23133\
        );

    \I__4646\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23133\
        );

    \I__4645\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23133\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__23147\,
            I => \N__23130\
        );

    \I__4643\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23127\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__23124\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__23130\,
            I => \N__23119\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__23127\,
            I => \N__23119\
        );

    \I__4639\ : Span4Mux_v
    port map (
            O => \N__23124\,
            I => \N__23116\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__23119\,
            I => \N__23113\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__23116\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__23113\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__23108\,
            I => \N__23100\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__23107\,
            I => \N__23096\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__23106\,
            I => \N__23093\
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__23105\,
            I => \N__23089\
        );

    \I__4631\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23078\
        );

    \I__4630\ : InMux
    port map (
            O => \N__23103\,
            I => \N__23078\
        );

    \I__4629\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23078\
        );

    \I__4628\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23078\
        );

    \I__4627\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23078\
        );

    \I__4626\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23071\
        );

    \I__4625\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23071\
        );

    \I__4624\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23071\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__23078\,
            I => \N__23066\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__23071\,
            I => \N__23066\
        );

    \I__4621\ : Span4Mux_h
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__23060\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1211\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__23057\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_0_cascade_\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_1_0_cascade_\
        );

    \I__4616\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__23048\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_0\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__23045\,
            I => \N__23042\
        );

    \I__4613\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__4611\ : Span4Mux_h
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__4610\ : Span4Mux_v
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__4609\ : Odrv4
    port map (
            O => \N__23030\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_0\
        );

    \I__4608\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23024\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__23024\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_0\
        );

    \I__4606\ : CascadeMux
    port map (
            O => \N__23021\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_0_cascade_\
        );

    \I__4605\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__23015\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_0\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__23012\,
            I => \N__23009\
        );

    \I__4602\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23006\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__23002\
        );

    \I__4600\ : InMux
    port map (
            O => \N__23005\,
            I => \N__22999\
        );

    \I__4599\ : Span4Mux_v
    port map (
            O => \N__23002\,
            I => \N__22996\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__22999\,
            I => \N__22993\
        );

    \I__4597\ : Span4Mux_s1_h
    port map (
            O => \N__22996\,
            I => \N__22990\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__22993\,
            I => \N__22987\
        );

    \I__4595\ : Span4Mux_h
    port map (
            O => \N__22990\,
            I => \N__22984\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__22987\,
            I => \processor_zipi8.sy_0\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__22984\,
            I => \processor_zipi8.sy_0\
        );

    \I__4592\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22975\
        );

    \I__4591\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22972\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__22975\,
            I => \N__22969\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__22972\,
            I => \N__22966\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__22969\,
            I => \N__22963\
        );

    \I__4587\ : Span4Mux_v
    port map (
            O => \N__22966\,
            I => \N__22960\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__22963\,
            I => \N__22957\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__22960\,
            I => \N__22954\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__22957\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__22954\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4\
        );

    \I__4582\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22945\
        );

    \I__4581\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22942\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__22945\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__22942\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5\
        );

    \I__4578\ : CEMux
    port map (
            O => \N__22937\,
            I => \N__22934\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__4576\ : Span4Mux_v
    port map (
            O => \N__22931\,
            I => \N__22927\
        );

    \I__4575\ : CEMux
    port map (
            O => \N__22930\,
            I => \N__22924\
        );

    \I__4574\ : Sp12to4
    port map (
            O => \N__22927\,
            I => \N__22921\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__22924\,
            I => \N__22918\
        );

    \I__4572\ : Odrv12
    port map (
            O => \N__22921\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__22918\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19\
        );

    \I__4570\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__22910\,
            I => \N__22906\
        );

    \I__4568\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22903\
        );

    \I__4567\ : Odrv12
    port map (
            O => \N__22906\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__22903\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6\
        );

    \I__4565\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22894\
        );

    \I__4564\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22891\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22888\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__22891\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6\
        );

    \I__4561\ : Odrv12
    port map (
            O => \N__22888\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__22883\,
            I => \N__22880\
        );

    \I__4559\ : InMux
    port map (
            O => \N__22880\,
            I => \N__22877\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__22877\,
            I => \N__22874\
        );

    \I__4557\ : Span12Mux_s3_h
    port map (
            O => \N__22874\,
            I => \N__22871\
        );

    \I__4556\ : Odrv12
    port map (
            O => \N__22871\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIUGIQ1_7\
        );

    \I__4555\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__22865\,
            I => \N__22862\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__4552\ : Odrv4
    port map (
            O => \N__22859\,
            I => \processor_zipi8.shift_rotate_result_7\
        );

    \I__4551\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22853\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__4549\ : Span4Mux_h
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__4548\ : Span4Mux_h
    port map (
            O => \N__22847\,
            I => \N__22844\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__22844\,
            I => \processor_zipi8.spm_data_7\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__22841\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269_cascade_\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__4544\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22829\
        );

    \I__4543\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22829\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__22829\,
            I => \N__22826\
        );

    \I__4541\ : Span4Mux_v
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__4540\ : Span4Mux_v
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__4539\ : Odrv4
    port map (
            O => \N__22820\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_7\
        );

    \I__4538\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22811\
        );

    \I__4537\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22811\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__22811\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_7\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__22808\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_243_cascade_\
        );

    \I__4534\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__4532\ : Span4Mux_h
    port map (
            O => \N__22799\,
            I => \N__22796\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__22796\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_299\
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__22793\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_5_cascade_\
        );

    \I__4529\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22787\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__4527\ : Span4Mux_s3_h
    port map (
            O => \N__22784\,
            I => \N__22781\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__4525\ : Span4Mux_v
    port map (
            O => \N__22778\,
            I => \N__22775\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__22775\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_315\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22765\
        );

    \I__4521\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22762\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__22765\,
            I => \N__22759\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22756\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__22759\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5\
        );

    \I__4517\ : Odrv12
    port map (
            O => \N__22756\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__22751\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_5_cascade_\
        );

    \I__4515\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22744\
        );

    \I__4514\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22741\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__22744\,
            I => \N__22736\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__22741\,
            I => \N__22736\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__22733\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_5\
        );

    \I__4509\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__22727\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_219\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__22724\,
            I => \N__22721\
        );

    \I__4506\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__22718\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_5\
        );

    \I__4504\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22712\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__22712\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_275\
        );

    \I__4502\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_5_cascade_\
        );

    \I__4501\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__22703\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_5\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_5_cascade_\
        );

    \I__4498\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__22694\,
            I => \N__22691\
        );

    \I__4496\ : Span4Mux_v
    port map (
            O => \N__22691\,
            I => \N__22688\
        );

    \I__4495\ : Span4Mux_h
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__22685\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_5\
        );

    \I__4493\ : InMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__22679\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_5\
        );

    \I__4491\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__22673\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_5\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__22670\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_5_cascade_\
        );

    \I__4488\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__22664\,
            I => \N__22660\
        );

    \I__4486\ : InMux
    port map (
            O => \N__22663\,
            I => \N__22657\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__22660\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__22657\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5\
        );

    \I__4483\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22649\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__22649\,
            I => \N__22645\
        );

    \I__4481\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22642\
        );

    \I__4480\ : Span4Mux_h
    port map (
            O => \N__22645\,
            I => \N__22637\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__22642\,
            I => \N__22637\
        );

    \I__4478\ : Span4Mux_v
    port map (
            O => \N__22637\,
            I => \N__22634\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__22634\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_5\
        );

    \I__4476\ : CascadeMux
    port map (
            O => \N__22631\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_5_cascade_\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__22628\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_6_cascade_\
        );

    \I__4474\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22622\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__22622\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI0VUU1_6\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__4471\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__4469\ : Span4Mux_v
    port map (
            O => \N__22610\,
            I => \N__22606\
        );

    \I__4468\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22603\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__22606\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__22603\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6\
        );

    \I__4465\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22595\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__22595\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIQCIQ1_6\
        );

    \I__4463\ : InMux
    port map (
            O => \N__22592\,
            I => \N__22588\
        );

    \I__4462\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22585\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__22588\,
            I => \N__22582\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__22585\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6\
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__22582\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6\
        );

    \I__4458\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22571\
        );

    \I__4457\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22571\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__22571\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_7\
        );

    \I__4455\ : SRMux
    port map (
            O => \N__22568\,
            I => \N__22564\
        );

    \I__4454\ : SRMux
    port map (
            O => \N__22567\,
            I => \N__22557\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__22564\,
            I => \N__22552\
        );

    \I__4452\ : SRMux
    port map (
            O => \N__22563\,
            I => \N__22549\
        );

    \I__4451\ : SRMux
    port map (
            O => \N__22562\,
            I => \N__22546\
        );

    \I__4450\ : SRMux
    port map (
            O => \N__22561\,
            I => \N__22543\
        );

    \I__4449\ : SRMux
    port map (
            O => \N__22560\,
            I => \N__22540\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__22557\,
            I => \N__22537\
        );

    \I__4447\ : SRMux
    port map (
            O => \N__22556\,
            I => \N__22534\
        );

    \I__4446\ : SRMux
    port map (
            O => \N__22555\,
            I => \N__22531\
        );

    \I__4445\ : Span4Mux_v
    port map (
            O => \N__22552\,
            I => \N__22524\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__22549\,
            I => \N__22524\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__22546\,
            I => \N__22521\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22516\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__22540\,
            I => \N__22516\
        );

    \I__4440\ : Span4Mux_s2_v
    port map (
            O => \N__22537\,
            I => \N__22509\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22509\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22509\
        );

    \I__4437\ : SRMux
    port map (
            O => \N__22530\,
            I => \N__22506\
        );

    \I__4436\ : SRMux
    port map (
            O => \N__22529\,
            I => \N__22503\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__22524\,
            I => \N__22498\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__22521\,
            I => \N__22493\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__22516\,
            I => \N__22493\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__22509\,
            I => \N__22486\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__22506\,
            I => \N__22486\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22486\
        );

    \I__4429\ : SRMux
    port map (
            O => \N__22502\,
            I => \N__22483\
        );

    \I__4428\ : SRMux
    port map (
            O => \N__22501\,
            I => \N__22480\
        );

    \I__4427\ : Span4Mux_v
    port map (
            O => \N__22498\,
            I => \N__22476\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__22493\,
            I => \N__22473\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__22486\,
            I => \N__22466\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22466\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__22480\,
            I => \N__22466\
        );

    \I__4422\ : SRMux
    port map (
            O => \N__22479\,
            I => \N__22463\
        );

    \I__4421\ : Sp12to4
    port map (
            O => \N__22476\,
            I => \N__22460\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__22473\,
            I => \N__22457\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__22466\,
            I => \N__22454\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__22463\,
            I => \N__22451\
        );

    \I__4417\ : Odrv12
    port map (
            O => \N__22460\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__22457\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__22454\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4414\ : Odrv12
    port map (
            O => \N__22451\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4413\ : InMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__22439\,
            I => \N__22435\
        );

    \I__4411\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22432\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__22435\,
            I => \N__22429\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__22432\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__22429\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__22424\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_6_cascade_\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNICIK32_6_cascade_\
        );

    \I__4405\ : CascadeMux
    port map (
            O => \N__22418\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_6_cascade_\
        );

    \I__4404\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__22406\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFJCI8_6\
        );

    \I__4400\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__22400\,
            I => \N__22396\
        );

    \I__4398\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22393\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__22396\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__22393\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2\
        );

    \I__4395\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22384\
        );

    \I__4394\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22381\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__22384\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__22381\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3\
        );

    \I__4391\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22372\
        );

    \I__4390\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22369\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__22372\,
            I => \N__22364\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__22369\,
            I => \N__22364\
        );

    \I__4387\ : Span4Mux_h
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__4386\ : Span4Mux_v
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__4385\ : Span4Mux_v
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__22355\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_6\
        );

    \I__4383\ : CEMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__4381\ : Span4Mux_s3_v
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__22340\,
            I => \N__22336\
        );

    \I__4378\ : CEMux
    port map (
            O => \N__22339\,
            I => \N__22333\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__22336\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__22333\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7\
        );

    \I__4375\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__4373\ : Span4Mux_h
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__4372\ : Span4Mux_v
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__22316\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI0ESR1_2\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__22313\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_2_cascade_\
        );

    \I__4369\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__22298\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI2HMP1_2\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__22295\,
            I => \N__22280\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__22294\,
            I => \N__22276\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__22293\,
            I => \N__22273\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__22292\,
            I => \N__22269\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__22291\,
            I => \N__22263\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__22290\,
            I => \N__22259\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__22289\,
            I => \N__22256\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__22288\,
            I => \N__22252\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__22287\,
            I => \N__22248\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__22286\,
            I => \N__22242\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__22285\,
            I => \N__22238\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__22284\,
            I => \N__22235\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__22283\,
            I => \N__22227\
        );

    \I__4351\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22210\
        );

    \I__4350\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22210\
        );

    \I__4349\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22210\
        );

    \I__4348\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22210\
        );

    \I__4347\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22210\
        );

    \I__4346\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22210\
        );

    \I__4345\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22210\
        );

    \I__4344\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22210\
        );

    \I__4343\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22193\
        );

    \I__4342\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22193\
        );

    \I__4341\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22193\
        );

    \I__4340\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22193\
        );

    \I__4339\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22193\
        );

    \I__4338\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22193\
        );

    \I__4337\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22193\
        );

    \I__4336\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22193\
        );

    \I__4335\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22176\
        );

    \I__4334\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22176\
        );

    \I__4333\ : InMux
    port map (
            O => \N__22246\,
            I => \N__22176\
        );

    \I__4332\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22176\
        );

    \I__4331\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22176\
        );

    \I__4330\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22176\
        );

    \I__4329\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22176\
        );

    \I__4328\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22176\
        );

    \I__4327\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22173\
        );

    \I__4326\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22170\
        );

    \I__4325\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22166\
        );

    \I__4324\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22163\
        );

    \I__4323\ : InMux
    port map (
            O => \N__22230\,
            I => \N__22160\
        );

    \I__4322\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22156\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__22210\,
            I => \N__22151\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__22193\,
            I => \N__22151\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__22176\,
            I => \N__22146\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__22173\,
            I => \N__22146\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__22170\,
            I => \N__22143\
        );

    \I__4316\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22140\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__22166\,
            I => \N__22129\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__22163\,
            I => \N__22124\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__22160\,
            I => \N__22124\
        );

    \I__4312\ : InMux
    port map (
            O => \N__22159\,
            I => \N__22121\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__22156\,
            I => \N__22116\
        );

    \I__4310\ : Sp12to4
    port map (
            O => \N__22151\,
            I => \N__22116\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__22146\,
            I => \N__22113\
        );

    \I__4308\ : Span4Mux_v
    port map (
            O => \N__22143\,
            I => \N__22110\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__22140\,
            I => \N__22107\
        );

    \I__4306\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22092\
        );

    \I__4305\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22092\
        );

    \I__4304\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22092\
        );

    \I__4303\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22092\
        );

    \I__4302\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22092\
        );

    \I__4301\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22092\
        );

    \I__4300\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22092\
        );

    \I__4299\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22089\
        );

    \I__4298\ : Span4Mux_s3_h
    port map (
            O => \N__22129\,
            I => \N__22082\
        );

    \I__4297\ : Span4Mux_v
    port map (
            O => \N__22124\,
            I => \N__22082\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22082\
        );

    \I__4295\ : Span12Mux_v
    port map (
            O => \N__22116\,
            I => \N__22079\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__22113\,
            I => \N__22076\
        );

    \I__4293\ : Span4Mux_v
    port map (
            O => \N__22110\,
            I => \N__22071\
        );

    \I__4292\ : Span4Mux_s3_v
    port map (
            O => \N__22107\,
            I => \N__22071\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22066\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22066\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__22082\,
            I => \N__22063\
        );

    \I__4288\ : Odrv12
    port map (
            O => \N__22079\,
            I => \processor_zipi8.sx_addr_4\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__22076\,
            I => \processor_zipi8.sx_addr_4\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__22071\,
            I => \processor_zipi8.sx_addr_4\
        );

    \I__4285\ : Odrv12
    port map (
            O => \N__22066\,
            I => \processor_zipi8.sx_addr_4\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__22063\,
            I => \processor_zipi8.sx_addr_4\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__22052\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI792G8_2_cascade_\
        );

    \I__4282\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__22046\,
            I => \N__22036\
        );

    \I__4280\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22031\
        );

    \I__4279\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22031\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__22043\,
            I => \N__22028\
        );

    \I__4277\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22019\
        );

    \I__4276\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22019\
        );

    \I__4275\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22019\
        );

    \I__4274\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22019\
        );

    \I__4273\ : Span4Mux_s3_h
    port map (
            O => \N__22036\,
            I => \N__22014\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__22031\,
            I => \N__22014\
        );

    \I__4271\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22010\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22007\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__22014\,
            I => \N__22004\
        );

    \I__4268\ : InMux
    port map (
            O => \N__22013\,
            I => \N__22001\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__21996\
        );

    \I__4266\ : Span4Mux_h
    port map (
            O => \N__22007\,
            I => \N__21996\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__22004\,
            I => \N__21993\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21990\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__21996\,
            I => \N__21987\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__21993\,
            I => \processor_zipi8.sx_2\
        );

    \I__4261\ : Odrv12
    port map (
            O => \N__21990\,
            I => \processor_zipi8.sx_2\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__21987\,
            I => \processor_zipi8.sx_2\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__21980\,
            I => \N__21976\
        );

    \I__4258\ : InMux
    port map (
            O => \N__21979\,
            I => \N__21973\
        );

    \I__4257\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21970\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__21973\,
            I => \N__21965\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__21970\,
            I => \N__21965\
        );

    \I__4254\ : Odrv12
    port map (
            O => \N__21965\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_0\
        );

    \I__4253\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__4251\ : Span12Mux_s8_h
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__4250\ : Odrv12
    port map (
            O => \N__21953\,
            I => \processor_zipi8.shift_rotate_result_3\
        );

    \I__4249\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__4247\ : Span4Mux_h
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__21938\,
            I => \processor_zipi8.spm_data_3\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__21935\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266_cascade_\
        );

    \I__4243\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21928\
        );

    \I__4242\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21925\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__21928\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__21925\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__4238\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__21914\,
            I => \N__21910\
        );

    \I__4236\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21907\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__21910\,
            I => \N__21902\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__21907\,
            I => \N__21902\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__21899\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_0\
        );

    \I__4231\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__21887\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI8MSR1_4\
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__4226\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21878\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__4224\ : Span4Mux_v
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__21872\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIAPMP1_4\
        );

    \I__4222\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__21866\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFIBI8_4\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__21863\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7A3G8_4_cascade_\
        );

    \I__4219\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21852\
        );

    \I__4217\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21847\
        );

    \I__4216\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21847\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__21852\,
            I => \N__21843\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21840\
        );

    \I__4213\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21837\
        );

    \I__4212\ : Span4Mux_s3_h
    port map (
            O => \N__21843\,
            I => \N__21828\
        );

    \I__4211\ : Span4Mux_v
    port map (
            O => \N__21840\,
            I => \N__21828\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__21837\,
            I => \N__21828\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__21836\,
            I => \N__21825\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__21835\,
            I => \N__21822\
        );

    \I__4207\ : Span4Mux_h
    port map (
            O => \N__21828\,
            I => \N__21818\
        );

    \I__4206\ : InMux
    port map (
            O => \N__21825\,
            I => \N__21811\
        );

    \I__4205\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21811\
        );

    \I__4204\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21811\
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__21818\,
            I => \processor_zipi8.sx_4\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__21811\,
            I => \processor_zipi8.sx_4\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__21806\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNISRE42_4_cascade_\
        );

    \I__4200\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__21800\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_4\
        );

    \I__4198\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__4196\ : Span4Mux_v
    port map (
            O => \N__21791\,
            I => \N__21787\
        );

    \I__4195\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21784\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__21787\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__21784\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__21779\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_2_cascade_\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__4190\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__21770\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_2\
        );

    \I__4188\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__4186\ : Odrv4
    port map (
            O => \N__21761\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI4KGN1_2\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__21758\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIKJE42_2_cascade_\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__21755\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_1_cascade_\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__21752\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_119_cascade_\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__21749\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_1_cascade_\
        );

    \I__4181\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__21743\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_95\
        );

    \I__4179\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__4177\ : Odrv12
    port map (
            O => \N__21734\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_151\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__4175\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__4173\ : Span4Mux_h
    port map (
            O => \N__21722\,
            I => \N__21719\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__21719\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_175\
        );

    \I__4171\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__21713\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_1\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__21710\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_191_cascade_\
        );

    \I__4168\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21703\
        );

    \I__4167\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21698\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__21703\,
            I => \N__21695\
        );

    \I__4165\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21690\
        );

    \I__4164\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21690\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__21698\,
            I => \N__21687\
        );

    \I__4162\ : Span4Mux_h
    port map (
            O => \N__21695\,
            I => \N__21677\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__21690\,
            I => \N__21677\
        );

    \I__4160\ : Span4Mux_v
    port map (
            O => \N__21687\,
            I => \N__21674\
        );

    \I__4159\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21669\
        );

    \I__4158\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21669\
        );

    \I__4157\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21662\
        );

    \I__4156\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21662\
        );

    \I__4155\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21662\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__21677\,
            I => \N__21655\
        );

    \I__4153\ : Span4Mux_h
    port map (
            O => \N__21674\,
            I => \N__21655\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__21669\,
            I => \N__21655\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__21662\,
            I => \processor_zipi8.sx_1\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__21655\,
            I => \processor_zipi8.sx_1\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__4148\ : InMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__4146\ : Odrv12
    port map (
            O => \N__21641\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNII4IQ1_4\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__4144\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__21629\,
            I => \N__21626\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__21626\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_4\
        );

    \I__4140\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__21620\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI4AK32_4\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__21617\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIOMUU1_4_cascade_\
        );

    \I__4137\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__21611\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_4\
        );

    \I__4135\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21604\
        );

    \I__4134\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21601\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__21604\,
            I => \N__21598\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__21601\,
            I => \N__21595\
        );

    \I__4131\ : Span4Mux_v
    port map (
            O => \N__21598\,
            I => \N__21592\
        );

    \I__4130\ : Odrv4
    port map (
            O => \N__21595\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__21592\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7\
        );

    \I__4128\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__21584\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_7\
        );

    \I__4126\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21575\
        );

    \I__4125\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21575\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__4123\ : Odrv12
    port map (
            O => \N__21572\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_7\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__21569\,
            I => \N__21566\
        );

    \I__4121\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21562\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__21565\,
            I => \N__21559\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21556\
        );

    \I__4118\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21553\
        );

    \I__4117\ : Span4Mux_v
    port map (
            O => \N__21556\,
            I => \N__21548\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__21553\,
            I => \N__21548\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__21548\,
            I => \N__21543\
        );

    \I__4114\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21538\
        );

    \I__4113\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21538\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__21543\,
            I => \processor_zipi8.port_id_1\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__21538\,
            I => \processor_zipi8.port_id_1\
        );

    \I__4110\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__4108\ : Span4Mux_h
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__21524\,
            I => \N__21521\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__21521\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_1\
        );

    \I__4105\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21509\
        );

    \I__4104\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21509\
        );

    \I__4103\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21509\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__21509\,
            I => \N__21504\
        );

    \I__4101\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21499\
        );

    \I__4100\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21499\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__21504\,
            I => \N__21494\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__21499\,
            I => \N__21494\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__4095\ : Span4Mux_s1_v
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__21485\,
            I => instruction_1
        );

    \I__4093\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__4091\ : Span4Mux_h
    port map (
            O => \N__21476\,
            I => \N__21473\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__21473\,
            I => \processor_zipi8.pc_vector_1\
        );

    \I__4089\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__21464\,
            I => \N__21461\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__21461\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_4\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__21458\,
            I => \N__21449\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__21457\,
            I => \N__21433\
        );

    \I__4083\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21429\
        );

    \I__4082\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21424\
        );

    \I__4081\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21424\
        );

    \I__4080\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21421\
        );

    \I__4079\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21418\
        );

    \I__4078\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21411\
        );

    \I__4077\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21411\
        );

    \I__4076\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21406\
        );

    \I__4075\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21406\
        );

    \I__4074\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21403\
        );

    \I__4073\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21392\
        );

    \I__4072\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21392\
        );

    \I__4071\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21392\
        );

    \I__4070\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21383\
        );

    \I__4069\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21383\
        );

    \I__4068\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21380\
        );

    \I__4067\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21375\
        );

    \I__4066\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21375\
        );

    \I__4065\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21372\
        );

    \I__4064\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21369\
        );

    \I__4063\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21366\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__21429\,
            I => \N__21357\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21357\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21357\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__21418\,
            I => \N__21357\
        );

    \I__4058\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21350\
        );

    \I__4057\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21350\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21345\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__21406\,
            I => \N__21345\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__21403\,
            I => \N__21342\
        );

    \I__4053\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21337\
        );

    \I__4052\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21337\
        );

    \I__4051\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21332\
        );

    \I__4050\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21332\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21329\
        );

    \I__4048\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21326\
        );

    \I__4047\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21319\
        );

    \I__4046\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21319\
        );

    \I__4045\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21319\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21316\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21311\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21311\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__21372\,
            I => \N__21306\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__21369\,
            I => \N__21306\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__21366\,
            I => \N__21301\
        );

    \I__4038\ : Span4Mux_v
    port map (
            O => \N__21357\,
            I => \N__21301\
        );

    \I__4037\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21296\
        );

    \I__4036\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21296\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__21350\,
            I => \N__21293\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__21345\,
            I => \N__21284\
        );

    \I__4033\ : Span4Mux_v
    port map (
            O => \N__21342\,
            I => \N__21284\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21284\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21284\
        );

    \I__4030\ : Span4Mux_s3_v
    port map (
            O => \N__21329\,
            I => \N__21281\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__21326\,
            I => \N__21274\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__21319\,
            I => \N__21274\
        );

    \I__4027\ : Span4Mux_h
    port map (
            O => \N__21316\,
            I => \N__21274\
        );

    \I__4026\ : Span4Mux_s3_v
    port map (
            O => \N__21311\,
            I => \N__21271\
        );

    \I__4025\ : Span4Mux_s3_v
    port map (
            O => \N__21306\,
            I => \N__21260\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__21301\,
            I => \N__21260\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__21296\,
            I => \N__21260\
        );

    \I__4022\ : Span4Mux_s3_v
    port map (
            O => \N__21293\,
            I => \N__21260\
        );

    \I__4021\ : Span4Mux_v
    port map (
            O => \N__21284\,
            I => \N__21260\
        );

    \I__4020\ : Span4Mux_h
    port map (
            O => \N__21281\,
            I => \N__21253\
        );

    \I__4019\ : Span4Mux_v
    port map (
            O => \N__21274\,
            I => \N__21253\
        );

    \I__4018\ : Span4Mux_h
    port map (
            O => \N__21271\,
            I => \N__21253\
        );

    \I__4017\ : Span4Mux_h
    port map (
            O => \N__21260\,
            I => \N__21250\
        );

    \I__4016\ : Odrv4
    port map (
            O => \N__21253\,
            I => instruction_12
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__21250\,
            I => instruction_12
        );

    \I__4014\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21239\
        );

    \I__4013\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21239\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__4010\ : Span4Mux_h
    port map (
            O => \N__21233\,
            I => \N__21230\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__21230\,
            I => \processor_zipi8.pc_vector_4\
        );

    \I__4008\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21220\
        );

    \I__4007\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21217\
        );

    \I__4006\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21204\
        );

    \I__4005\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21204\
        );

    \I__4004\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21204\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__21220\,
            I => \N__21201\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__21217\,
            I => \N__21198\
        );

    \I__4001\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21193\
        );

    \I__4000\ : InMux
    port map (
            O => \N__21215\,
            I => \N__21193\
        );

    \I__3999\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21190\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__21213\,
            I => \N__21186\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__21212\,
            I => \N__21183\
        );

    \I__3996\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21176\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__21204\,
            I => \N__21171\
        );

    \I__3994\ : Span4Mux_v
    port map (
            O => \N__21201\,
            I => \N__21171\
        );

    \I__3993\ : Span4Mux_h
    port map (
            O => \N__21198\,
            I => \N__21164\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__21193\,
            I => \N__21164\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__21190\,
            I => \N__21164\
        );

    \I__3990\ : InMux
    port map (
            O => \N__21189\,
            I => \N__21157\
        );

    \I__3989\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21157\
        );

    \I__3988\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21157\
        );

    \I__3987\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21152\
        );

    \I__3986\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21152\
        );

    \I__3985\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21147\
        );

    \I__3984\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21147\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__21176\,
            I => \N__21144\
        );

    \I__3982\ : Span4Mux_v
    port map (
            O => \N__21171\,
            I => \N__21135\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__21164\,
            I => \N__21135\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__21157\,
            I => \N__21135\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N__21135\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__21147\,
            I => \N__21132\
        );

    \I__3977\ : Span4Mux_s2_v
    port map (
            O => \N__21144\,
            I => \N__21129\
        );

    \I__3976\ : Span4Mux_s2_v
    port map (
            O => \N__21135\,
            I => \N__21124\
        );

    \I__3975\ : Span4Mux_h
    port map (
            O => \N__21132\,
            I => \N__21124\
        );

    \I__3974\ : Span4Mux_h
    port map (
            O => \N__21129\,
            I => \N__21121\
        );

    \I__3973\ : Span4Mux_h
    port map (
            O => \N__21124\,
            I => \N__21118\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__21121\,
            I => instruction_13
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__21118\,
            I => instruction_13
        );

    \I__3970\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21107\
        );

    \I__3969\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21103\
        );

    \I__3968\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21100\
        );

    \I__3967\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21097\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__21107\,
            I => \N__21094\
        );

    \I__3965\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21091\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__21103\,
            I => \N__21087\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__21100\,
            I => \N__21084\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__21097\,
            I => \N__21075\
        );

    \I__3961\ : Span4Mux_s3_h
    port map (
            O => \N__21094\,
            I => \N__21072\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__21091\,
            I => \N__21069\
        );

    \I__3959\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21066\
        );

    \I__3958\ : Span4Mux_v
    port map (
            O => \N__21087\,
            I => \N__21061\
        );

    \I__3957\ : Span4Mux_s3_h
    port map (
            O => \N__21084\,
            I => \N__21061\
        );

    \I__3956\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21058\
        );

    \I__3955\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21047\
        );

    \I__3954\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21047\
        );

    \I__3953\ : InMux
    port map (
            O => \N__21080\,
            I => \N__21047\
        );

    \I__3952\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21047\
        );

    \I__3951\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21047\
        );

    \I__3950\ : Odrv12
    port map (
            O => \N__21075\,
            I => \processor_zipi8.sx_0\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__21072\,
            I => \processor_zipi8.sx_0\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__21069\,
            I => \processor_zipi8.sx_0\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__21066\,
            I => \processor_zipi8.sx_0\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__21061\,
            I => \processor_zipi8.sx_0\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__21058\,
            I => \processor_zipi8.sx_0\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__21047\,
            I => \processor_zipi8.sx_0\
        );

    \I__3943\ : IoInMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__3941\ : IoSpan4Mux
    port map (
            O => \N__21026\,
            I => \N__21023\
        );

    \I__3940\ : Span4Mux_s3_h
    port map (
            O => \N__21023\,
            I => \N__21020\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__21020\,
            I => \LED1_c\
        );

    \I__3938\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21011\
        );

    \I__3937\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21011\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__3935\ : Span12Mux_s10_h
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__3934\ : Odrv12
    port map (
            O => \N__21005\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_1\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__21002\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_1_cascade_\
        );

    \I__3932\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20993\
        );

    \I__3931\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20993\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__3929\ : Odrv12
    port map (
            O => \N__20990\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_1\
        );

    \I__3928\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__20984\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1\
        );

    \I__3926\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20975\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20975\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__20972\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_1\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__3921\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20960\
        );

    \I__3920\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20960\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__20960\,
            I => \N__20957\
        );

    \I__3918\ : Span4Mux_v
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__20954\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_1\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__20951\,
            I => \N__20948\
        );

    \I__3915\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__20945\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_1\
        );

    \I__3913\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__3911\ : Odrv12
    port map (
            O => \N__20936\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_7\
        );

    \I__3910\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20930\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__3908\ : Span4Mux_s3_h
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__20921\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_7\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__20918\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_0_cascade_\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__20915\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_0_cascade_\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__3902\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__20906\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_7\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__20903\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_0_cascade_\
        );

    \I__3899\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__20897\,
            I => \N__20893\
        );

    \I__3897\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__20893\,
            I => \N__20885\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__20890\,
            I => \N__20885\
        );

    \I__3894\ : Span4Mux_v
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__20882\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_0\
        );

    \I__3892\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__20876\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_0\
        );

    \I__3890\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20867\
        );

    \I__3889\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20867\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__3887\ : Span4Mux_h
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__20861\,
            I => \processor_zipi8.register_enable\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__20858\,
            I => \N__20843\
        );

    \I__3884\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20832\
        );

    \I__3883\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20832\
        );

    \I__3882\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20832\
        );

    \I__3881\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20832\
        );

    \I__3880\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20828\
        );

    \I__3879\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20813\
        );

    \I__3878\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20813\
        );

    \I__3877\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20813\
        );

    \I__3876\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20813\
        );

    \I__3875\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20813\
        );

    \I__3874\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20813\
        );

    \I__3873\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20813\
        );

    \I__3872\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20808\
        );

    \I__3871\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20808\
        );

    \I__3870\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20805\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__20832\,
            I => \N__20802\
        );

    \I__3868\ : InMux
    port map (
            O => \N__20831\,
            I => \N__20799\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__20828\,
            I => \N__20794\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__20813\,
            I => \N__20794\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__20808\,
            I => \N__20787\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20787\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__20802\,
            I => \N__20787\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20782\
        );

    \I__3861\ : Sp12to4
    port map (
            O => \N__20794\,
            I => \N__20782\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__20787\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205\
        );

    \I__3859\ : Odrv12
    port map (
            O => \N__20782\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205\
        );

    \I__3858\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__20771\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_0\
        );

    \I__3855\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__20765\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNISBGN1_0\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__20762\,
            I => \N__20759\
        );

    \I__3852\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__20756\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_1\
        );

    \I__3850\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20749\
        );

    \I__3849\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20746\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20740\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__20743\,
            I => \N__20735\
        );

    \I__3845\ : Span4Mux_h
    port map (
            O => \N__20740\,
            I => \N__20735\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__20735\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_1\
        );

    \I__3843\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20728\
        );

    \I__3842\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20725\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__20728\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__20725\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1\
        );

    \I__3839\ : CascadeMux
    port map (
            O => \N__20720\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_1_cascade_\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__20717\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_cascade_\
        );

    \I__3837\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20708\
        );

    \I__3836\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20708\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__3834\ : Span4Mux_v
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__3833\ : Span4Mux_h
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__20699\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_1\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__20696\,
            I => \N__20692\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__20695\,
            I => \N__20689\
        );

    \I__3829\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20684\
        );

    \I__3828\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20684\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__20684\,
            I => \N__20681\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__20678\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_1\
        );

    \I__3824\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__20672\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_5\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__20669\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_5_cascade_\
        );

    \I__3821\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20663\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__20663\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_5\
        );

    \I__3819\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20648\
        );

    \I__3818\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20648\
        );

    \I__3817\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20648\
        );

    \I__3816\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20648\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__20648\,
            I => \N__20635\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__20647\,
            I => \N__20632\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__20646\,
            I => \N__20629\
        );

    \I__3812\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20624\
        );

    \I__3811\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20609\
        );

    \I__3810\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20609\
        );

    \I__3809\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20609\
        );

    \I__3808\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20609\
        );

    \I__3807\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20609\
        );

    \I__3806\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20609\
        );

    \I__3805\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20609\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__20635\,
            I => \N__20606\
        );

    \I__3803\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20597\
        );

    \I__3802\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20597\
        );

    \I__3801\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20597\
        );

    \I__3800\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20597\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__20624\,
            I => \N__20592\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20592\
        );

    \I__3797\ : Sp12to4
    port map (
            O => \N__20606\,
            I => \N__20587\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__20597\,
            I => \N__20587\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__20592\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206\
        );

    \I__3794\ : Odrv12
    port map (
            O => \N__20587\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206\
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__20582\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_0_cascade_\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__20579\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNICBE42_0_cascade_\
        );

    \I__3791\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20570\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__20567\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIQ8MP1_0\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__20564\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_0_cascade_\
        );

    \I__3786\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__20558\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIO5SR1_0\
        );

    \I__3784\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__20546\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI781G8_0\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__20543\,
            I => \N__20536\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__20542\,
            I => \N__20531\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__20541\,
            I => \N__20528\
        );

    \I__3777\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20524\
        );

    \I__3776\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20519\
        );

    \I__3775\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20519\
        );

    \I__3774\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20514\
        );

    \I__3773\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20514\
        );

    \I__3772\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20507\
        );

    \I__3771\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20507\
        );

    \I__3770\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20507\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__20524\,
            I => \N__20502\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20502\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20497\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__20507\,
            I => \N__20497\
        );

    \I__3765\ : Span4Mux_v
    port map (
            O => \N__20502\,
            I => \N__20494\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__20497\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__20494\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209\
        );

    \I__3762\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20486\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20482\
        );

    \I__3760\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20479\
        );

    \I__3759\ : Span4Mux_h
    port map (
            O => \N__20482\,
            I => \N__20474\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__20479\,
            I => \N__20474\
        );

    \I__3757\ : Span4Mux_v
    port map (
            O => \N__20474\,
            I => \N__20471\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__20471\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_7\
        );

    \I__3755\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20462\
        );

    \I__3754\ : InMux
    port map (
            O => \N__20467\,
            I => \N__20462\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__20459\,
            I => \N__20456\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__20456\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_7\
        );

    \I__3750\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20450\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__3748\ : Span4Mux_s3_h
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__20444\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_7\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__20441\,
            I => \N__20437\
        );

    \I__3745\ : InMux
    port map (
            O => \N__20440\,
            I => \N__20432\
        );

    \I__3744\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20432\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__20429\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_7\
        );

    \I__3741\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20420\
        );

    \I__3740\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20420\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__3738\ : Span4Mux_v
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__20414\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_7\
        );

    \I__3736\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__3734\ : Odrv12
    port map (
            O => \N__20405\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_7\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__20402\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_5_cascade_\
        );

    \I__3732\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__3730\ : Span12Mux_s6_h
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__3729\ : Odrv12
    port map (
            O => \N__20390\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_5\
        );

    \I__3728\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20383\
        );

    \I__3727\ : InMux
    port map (
            O => \N__20386\,
            I => \N__20380\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__20383\,
            I => \N__20377\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__20380\,
            I => \N__20372\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__20377\,
            I => \N__20372\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__20372\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_0\
        );

    \I__3722\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20365\
        );

    \I__3721\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20362\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__20365\,
            I => \N__20359\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__20362\,
            I => \N__20356\
        );

    \I__3718\ : Span4Mux_h
    port map (
            O => \N__20359\,
            I => \N__20351\
        );

    \I__3717\ : Span4Mux_v
    port map (
            O => \N__20356\,
            I => \N__20351\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__20351\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_0\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__3714\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__20342\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_0\
        );

    \I__3712\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__20336\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_5\
        );

    \I__3710\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20327\
        );

    \I__3709\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20327\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20321\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__20326\,
            I => \N__20318\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N__20313\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \N__20310\
        );

    \I__3704\ : Span4Mux_h
    port map (
            O => \N__20321\,
            I => \N__20307\
        );

    \I__3703\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20304\
        );

    \I__3702\ : InMux
    port map (
            O => \N__20317\,
            I => \N__20295\
        );

    \I__3701\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20295\
        );

    \I__3700\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20295\
        );

    \I__3699\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20295\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__20307\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__20304\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__20295\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212\
        );

    \I__3695\ : CEMux
    port map (
            O => \N__20288\,
            I => \N__20284\
        );

    \I__3694\ : CEMux
    port map (
            O => \N__20287\,
            I => \N__20281\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__20284\,
            I => \N__20278\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20275\
        );

    \I__3691\ : Span4Mux_v
    port map (
            O => \N__20278\,
            I => \N__20272\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__20275\,
            I => \N__20269\
        );

    \I__3689\ : Span4Mux_h
    port map (
            O => \N__20272\,
            I => \N__20266\
        );

    \I__3688\ : Span4Mux_h
    port map (
            O => \N__20269\,
            I => \N__20263\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__20266\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__20263\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__20258\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_4_cascade_\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__20255\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_7_cascade_\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__3682\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20246\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__3680\ : Span12Mux_s6_h
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__3679\ : Odrv12
    port map (
            O => \N__20240\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIO8HN1_7\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__20237\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_7_cascade_\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__20234\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_7_cascade_\
        );

    \I__3676\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__20228\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI43VU1_7\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__20225\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIGMK32_7_cascade_\
        );

    \I__3673\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__3671\ : Span4Mux_v
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__3670\ : Span4Mux_h
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__20207\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_7\
        );

    \I__3667\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20200\
        );

    \I__3666\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20197\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__20200\,
            I => \N__20194\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__20197\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__20194\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__20189\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_7_cascade_\
        );

    \I__3661\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20180\
        );

    \I__3660\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20180\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__3658\ : Span4Mux_h
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__20174\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_7\
        );

    \I__3656\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20168\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__20168\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_7\
        );

    \I__3654\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20161\
        );

    \I__3653\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20158\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__20161\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__20158\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__3649\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__20144\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_3\
        );

    \I__3646\ : CEMux
    port map (
            O => \N__20141\,
            I => \N__20137\
        );

    \I__3645\ : CEMux
    port map (
            O => \N__20140\,
            I => \N__20134\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N__20131\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20128\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__20131\,
            I => \N__20125\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__20128\,
            I => \N__20122\
        );

    \I__3640\ : Span4Mux_s1_v
    port map (
            O => \N__20125\,
            I => \N__20119\
        );

    \I__3639\ : Span4Mux_v
    port map (
            O => \N__20122\,
            I => \N__20116\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__20119\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__20116\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6\
        );

    \I__3636\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__20108\,
            I => \processor_zipi8.alu_result_4\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__20105\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI8OGN1_3_cascade_\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__20102\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_am_1_3_cascade_\
        );

    \I__3632\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__20096\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIONE42_3\
        );

    \I__3630\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__20090\,
            I => \N__20087\
        );

    \I__3628\ : Span12Mux_s3_v
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__3627\ : Odrv12
    port map (
            O => \N__20084\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI6LMP1_3\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__3625\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__3623\ : Span12Mux_s5_v
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__3622\ : Odrv12
    port map (
            O => \N__20069\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI4ISR1_3\
        );

    \I__3621\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__20063\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_3\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__20060\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINP2G8_3_cascade_\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__20057\,
            I => \N__20053\
        );

    \I__3617\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20047\
        );

    \I__3616\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20040\
        );

    \I__3615\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20040\
        );

    \I__3614\ : InMux
    port map (
            O => \N__20051\,
            I => \N__20037\
        );

    \I__3613\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20034\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__20047\,
            I => \N__20031\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__20046\,
            I => \N__20028\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__20045\,
            I => \N__20025\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__20021\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__20018\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20015\
        );

    \I__3606\ : Span4Mux_h
    port map (
            O => \N__20031\,
            I => \N__20011\
        );

    \I__3605\ : InMux
    port map (
            O => \N__20028\,
            I => \N__20004\
        );

    \I__3604\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20004\
        );

    \I__3603\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20004\
        );

    \I__3602\ : Span12Mux_s5_h
    port map (
            O => \N__20021\,
            I => \N__20001\
        );

    \I__3601\ : Span4Mux_h
    port map (
            O => \N__20018\,
            I => \N__19996\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__20015\,
            I => \N__19996\
        );

    \I__3599\ : InMux
    port map (
            O => \N__20014\,
            I => \N__19993\
        );

    \I__3598\ : Span4Mux_v
    port map (
            O => \N__20011\,
            I => \N__19988\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__19988\
        );

    \I__3596\ : Odrv12
    port map (
            O => \N__20001\,
            I => \processor_zipi8.sx_3\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__19996\,
            I => \processor_zipi8.sx_3\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__19993\,
            I => \processor_zipi8.sx_3\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__19988\,
            I => \processor_zipi8.sx_3\
        );

    \I__3592\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__3590\ : Odrv12
    port map (
            O => \N__19973\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_4\
        );

    \I__3589\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__19967\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_4\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19960\
        );

    \I__3586\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19955\
        );

    \I__3585\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19952\
        );

    \I__3584\ : CascadeMux
    port map (
            O => \N__19959\,
            I => \N__19940\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \N__19933\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__19955\,
            I => \N__19926\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19926\
        );

    \I__3580\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19919\
        );

    \I__3579\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19919\
        );

    \I__3578\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19919\
        );

    \I__3577\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19914\
        );

    \I__3576\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19909\
        );

    \I__3575\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19909\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19904\
        );

    \I__3573\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19904\
        );

    \I__3572\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19898\
        );

    \I__3571\ : InMux
    port map (
            O => \N__19940\,
            I => \N__19887\
        );

    \I__3570\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19887\
        );

    \I__3569\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19887\
        );

    \I__3568\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19887\
        );

    \I__3567\ : InMux
    port map (
            O => \N__19936\,
            I => \N__19887\
        );

    \I__3566\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19880\
        );

    \I__3565\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19880\
        );

    \I__3564\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19880\
        );

    \I__3563\ : Span4Mux_v
    port map (
            O => \N__19926\,
            I => \N__19875\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19875\
        );

    \I__3561\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19872\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__19917\,
            I => \N__19866\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__19914\,
            I => \N__19859\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19859\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19859\
        );

    \I__3556\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19852\
        );

    \I__3555\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19852\
        );

    \I__3554\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19852\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19845\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__19887\,
            I => \N__19845\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19845\
        );

    \I__3550\ : Span4Mux_h
    port map (
            O => \N__19875\,
            I => \N__19842\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__19872\,
            I => \N__19839\
        );

    \I__3548\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19830\
        );

    \I__3547\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19830\
        );

    \I__3546\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19830\
        );

    \I__3545\ : InMux
    port map (
            O => \N__19866\,
            I => \N__19830\
        );

    \I__3544\ : Span4Mux_v
    port map (
            O => \N__19859\,
            I => \N__19827\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__19852\,
            I => \N__19824\
        );

    \I__3542\ : Span4Mux_h
    port map (
            O => \N__19845\,
            I => \N__19819\
        );

    \I__3541\ : Span4Mux_v
    port map (
            O => \N__19842\,
            I => \N__19819\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__19839\,
            I => \N__19816\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__19830\,
            I => \N__19809\
        );

    \I__3538\ : Sp12to4
    port map (
            O => \N__19827\,
            I => \N__19809\
        );

    \I__3537\ : Span12Mux_s2_h
    port map (
            O => \N__19824\,
            I => \N__19809\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__19819\,
            I => \N__19806\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__19816\,
            I => instruction_14
        );

    \I__3534\ : Odrv12
    port map (
            O => \N__19809\,
            I => instruction_14
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__19806\,
            I => instruction_14
        );

    \I__3532\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19791\
        );

    \I__3531\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19788\
        );

    \I__3530\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19785\
        );

    \I__3529\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19771\
        );

    \I__3528\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19771\
        );

    \I__3527\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19768\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__19791\,
            I => \N__19761\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__19788\,
            I => \N__19761\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19761\
        );

    \I__3523\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19758\
        );

    \I__3522\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19755\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__19782\,
            I => \N__19752\
        );

    \I__3520\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19744\
        );

    \I__3519\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19744\
        );

    \I__3518\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19744\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__19778\,
            I => \N__19740\
        );

    \I__3516\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19734\
        );

    \I__3515\ : InMux
    port map (
            O => \N__19776\,
            I => \N__19734\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19729\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__19768\,
            I => \N__19729\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__19761\,
            I => \N__19722\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__19758\,
            I => \N__19722\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19722\
        );

    \I__3509\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19717\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19717\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19714\
        );

    \I__3506\ : InMux
    port map (
            O => \N__19743\,
            I => \N__19709\
        );

    \I__3505\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19709\
        );

    \I__3504\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19706\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__19734\,
            I => \N__19701\
        );

    \I__3502\ : Span4Mux_h
    port map (
            O => \N__19729\,
            I => \N__19701\
        );

    \I__3501\ : Span4Mux_h
    port map (
            O => \N__19722\,
            I => \N__19698\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19691\
        );

    \I__3499\ : Span4Mux_h
    port map (
            O => \N__19714\,
            I => \N__19691\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__19709\,
            I => \N__19691\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__19706\,
            I => \processor_zipi8.arith_logical_sel_1_0_2\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__19701\,
            I => \processor_zipi8.arith_logical_sel_1_0_2\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__19698\,
            I => \processor_zipi8.arith_logical_sel_1_0_2\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__19691\,
            I => \processor_zipi8.arith_logical_sel_1_0_2\
        );

    \I__3493\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__3491\ : Span12Mux_s6_v
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__3490\ : Odrv12
    port map (
            O => \N__19673\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_3\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__19670\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_3_cascade_\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__19667\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_3_cascade_\
        );

    \I__3487\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__19661\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_3\
        );

    \I__3485\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__19655\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_3\
        );

    \I__3483\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19646\
        );

    \I__3482\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19646\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__19646\,
            I => \processor_zipi8.sy_3\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__19643\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_bm_1_3_cascade_\
        );

    \I__3479\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19636\
        );

    \I__3478\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19633\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__19636\,
            I => \N__19628\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__19633\,
            I => \N__19625\
        );

    \I__3475\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19622\
        );

    \I__3474\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19619\
        );

    \I__3473\ : Span4Mux_v
    port map (
            O => \N__19628\,
            I => \N__19614\
        );

    \I__3472\ : Span12Mux_s9_v
    port map (
            O => \N__19625\,
            I => \N__19609\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__19622\,
            I => \N__19609\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__19619\,
            I => \N__19606\
        );

    \I__3469\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19603\
        );

    \I__3468\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19600\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__19614\,
            I => \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical\
        );

    \I__3466\ : Odrv12
    port map (
            O => \N__19609\,
            I => \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical\
        );

    \I__3465\ : Odrv12
    port map (
            O => \N__19606\,
            I => \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__19603\,
            I => \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__19600\,
            I => \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical\
        );

    \I__3462\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19581\
        );

    \I__3461\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19581\
        );

    \I__3460\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19572\
        );

    \I__3459\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19572\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__19581\,
            I => \N__19569\
        );

    \I__3457\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19564\
        );

    \I__3456\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19564\
        );

    \I__3455\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19558\
        );

    \I__3454\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19558\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__19572\,
            I => \N__19552\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__19569\,
            I => \N__19546\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__19564\,
            I => \N__19546\
        );

    \I__3450\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19543\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19540\
        );

    \I__3448\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19537\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__19556\,
            I => \N__19533\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__19555\,
            I => \N__19530\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__19552\,
            I => \N__19527\
        );

    \I__3444\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19524\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__19546\,
            I => \N__19515\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__19543\,
            I => \N__19515\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__19540\,
            I => \N__19515\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__19537\,
            I => \N__19515\
        );

    \I__3439\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19508\
        );

    \I__3438\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19508\
        );

    \I__3437\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19508\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__19527\,
            I => \processor_zipi8.un4_arith_logical_sel\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__19524\,
            I => \processor_zipi8.un4_arith_logical_sel\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__19515\,
            I => \processor_zipi8.un4_arith_logical_sel\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__19508\,
            I => \processor_zipi8.un4_arith_logical_sel\
        );

    \I__3432\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__19496\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1Z0Z_1\
        );

    \I__3430\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__19490\,
            I => \processor_zipi8.arith_and_logic_operations_i.N_773_tz\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__19487\,
            I => \N__19483\
        );

    \I__3427\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19479\
        );

    \I__3426\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19475\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__19482\,
            I => \N__19468\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__19479\,
            I => \N__19464\
        );

    \I__3423\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19461\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__19475\,
            I => \N__19458\
        );

    \I__3421\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19454\
        );

    \I__3420\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19451\
        );

    \I__3419\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19444\
        );

    \I__3418\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19444\
        );

    \I__3417\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19444\
        );

    \I__3416\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19441\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__19464\,
            I => \N__19434\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__19461\,
            I => \N__19434\
        );

    \I__3413\ : Span4Mux_v
    port map (
            O => \N__19458\,
            I => \N__19434\
        );

    \I__3412\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19431\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__19454\,
            I => \N__19428\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__19451\,
            I => \N__19425\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__19444\,
            I => \N__19420\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__19441\,
            I => \N__19420\
        );

    \I__3407\ : Span4Mux_h
    port map (
            O => \N__19434\,
            I => \N__19415\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__19431\,
            I => \N__19415\
        );

    \I__3405\ : Span12Mux_v
    port map (
            O => \N__19428\,
            I => \N__19412\
        );

    \I__3404\ : Span4Mux_v
    port map (
            O => \N__19425\,
            I => \N__19407\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__19420\,
            I => \N__19407\
        );

    \I__3402\ : Span4Mux_v
    port map (
            O => \N__19415\,
            I => \N__19404\
        );

    \I__3401\ : Odrv12
    port map (
            O => \N__19412\,
            I => \processor_zipi8.arith_logical_sel_1_0_0\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__19407\,
            I => \processor_zipi8.arith_logical_sel_1_0_0\
        );

    \I__3399\ : Odrv4
    port map (
            O => \N__19404\,
            I => \processor_zipi8.arith_logical_sel_1_0_0\
        );

    \I__3398\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__19394\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_1\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__19391\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_4_cascade_\
        );

    \I__3395\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__19382\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_4\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__19379\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_4_cascade_\
        );

    \I__3391\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19370\
        );

    \I__3390\ : InMux
    port map (
            O => \N__19375\,
            I => \N__19370\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__3388\ : Span4Mux_v
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__19361\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_4\
        );

    \I__3385\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__19355\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_4\
        );

    \I__3383\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__19349\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_4\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__19346\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_4_cascade_\
        );

    \I__3380\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__19337\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_4\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__19334\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4_cascade_\
        );

    \I__3376\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19325\
        );

    \I__3375\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19325\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__19325\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_34_5\
        );

    \I__3373\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19316\
        );

    \I__3372\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19316\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__3370\ : Odrv12
    port map (
            O => \N__19313\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_5\
        );

    \I__3369\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__19307\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4\
        );

    \I__3367\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__19301\,
            I => \processor_zipi8.flags_i.parity_5\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__19298\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_1_cascade_\
        );

    \I__3364\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19291\
        );

    \I__3363\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19288\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__19291\,
            I => \processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__19288\,
            I => \processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1\
        );

    \I__3360\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__19280\,
            I => \N__19276\
        );

    \I__3358\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19273\
        );

    \I__3357\ : Odrv12
    port map (
            O => \N__19276\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__19273\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1\
        );

    \I__3355\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__19265\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tzZ0Z_4\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__19262\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_4_cascade_\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__19259\,
            I => \N__19255\
        );

    \I__3351\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19250\
        );

    \I__3350\ : InMux
    port map (
            O => \N__19255\,
            I => \N__19250\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__19250\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_4\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__19247\,
            I => \N__19243\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__19246\,
            I => \N__19240\
        );

    \I__3346\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19237\
        );

    \I__3345\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19231\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__19237\,
            I => \N__19228\
        );

    \I__3343\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19221\
        );

    \I__3342\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19221\
        );

    \I__3341\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19221\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__19231\,
            I => \N__19218\
        );

    \I__3339\ : Span4Mux_h
    port map (
            O => \N__19228\,
            I => \N__19213\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__19221\,
            I => \N__19213\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__19218\,
            I => \processor_zipi8.port_id_4\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__19213\,
            I => \processor_zipi8.port_id_4\
        );

    \I__3335\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19195\
        );

    \I__3334\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19195\
        );

    \I__3333\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19190\
        );

    \I__3332\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19190\
        );

    \I__3331\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19181\
        );

    \I__3330\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19181\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__19202\,
            I => \N__19177\
        );

    \I__3328\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19172\
        );

    \I__3327\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19172\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__19195\,
            I => \N__19167\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__19190\,
            I => \N__19167\
        );

    \I__3324\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19160\
        );

    \I__3323\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19160\
        );

    \I__3322\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19160\
        );

    \I__3321\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19157\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__19181\,
            I => \N__19154\
        );

    \I__3319\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19147\
        );

    \I__3318\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19147\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__19172\,
            I => \N__19144\
        );

    \I__3316\ : Span4Mux_h
    port map (
            O => \N__19167\,
            I => \N__19137\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__19160\,
            I => \N__19137\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__19157\,
            I => \N__19137\
        );

    \I__3313\ : Span4Mux_v
    port map (
            O => \N__19154\,
            I => \N__19134\
        );

    \I__3312\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19129\
        );

    \I__3311\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19129\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__19147\,
            I => \N__19126\
        );

    \I__3309\ : Span4Mux_v
    port map (
            O => \N__19144\,
            I => \N__19121\
        );

    \I__3308\ : Span4Mux_v
    port map (
            O => \N__19137\,
            I => \N__19121\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__19134\,
            I => \processor_zipi8.arith_logical_sel_1\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__19129\,
            I => \processor_zipi8.arith_logical_sel_1\
        );

    \I__3305\ : Odrv12
    port map (
            O => \N__19126\,
            I => \processor_zipi8.arith_logical_sel_1\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__19121\,
            I => \processor_zipi8.arith_logical_sel_1\
        );

    \I__3303\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__19109\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_4\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__19106\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198_cascade_\
        );

    \I__3300\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19099\
        );

    \I__3299\ : InMux
    port map (
            O => \N__19102\,
            I => \N__19096\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__19099\,
            I => \N__19093\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__19096\,
            I => \N__19090\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__19093\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__19090\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3\
        );

    \I__3294\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__19082\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__3291\ : InMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__19073\,
            I => \processor_zipi8.decode4_strobes_enables_i.un8_register_enable_type\
        );

    \I__3289\ : CEMux
    port map (
            O => \N__19070\,
            I => \N__19062\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \N__19053\
        );

    \I__3287\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19046\
        );

    \I__3286\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19046\
        );

    \I__3285\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19046\
        );

    \I__3284\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19043\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__19062\,
            I => \N__19038\
        );

    \I__3282\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19035\
        );

    \I__3281\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19032\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__19059\,
            I => \N__19028\
        );

    \I__3279\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19025\
        );

    \I__3278\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19018\
        );

    \I__3277\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19018\
        );

    \I__3276\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19018\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__19046\,
            I => \N__19013\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__19043\,
            I => \N__19013\
        );

    \I__3273\ : InMux
    port map (
            O => \N__19042\,
            I => \N__19010\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__19041\,
            I => \N__19006\
        );

    \I__3271\ : Span4Mux_v
    port map (
            O => \N__19038\,
            I => \N__19002\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__19035\,
            I => \N__18995\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__19032\,
            I => \N__18995\
        );

    \I__3268\ : InMux
    port map (
            O => \N__19031\,
            I => \N__18992\
        );

    \I__3267\ : InMux
    port map (
            O => \N__19028\,
            I => \N__18989\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__19025\,
            I => \N__18980\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__19018\,
            I => \N__18980\
        );

    \I__3264\ : Span4Mux_h
    port map (
            O => \N__19013\,
            I => \N__18980\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__19010\,
            I => \N__18980\
        );

    \I__3262\ : InMux
    port map (
            O => \N__19009\,
            I => \N__18977\
        );

    \I__3261\ : InMux
    port map (
            O => \N__19006\,
            I => \N__18972\
        );

    \I__3260\ : InMux
    port map (
            O => \N__19005\,
            I => \N__18972\
        );

    \I__3259\ : Span4Mux_s2_h
    port map (
            O => \N__19002\,
            I => \N__18969\
        );

    \I__3258\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18964\
        );

    \I__3257\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18964\
        );

    \I__3256\ : Span4Mux_v
    port map (
            O => \N__18995\,
            I => \N__18961\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__18992\,
            I => \N__18956\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__18989\,
            I => \N__18956\
        );

    \I__3253\ : Span4Mux_v
    port map (
            O => \N__18980\,
            I => \N__18953\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__18977\,
            I => \N__18950\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__18972\,
            I => \processor_zipi8.t_state_1\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__18969\,
            I => \processor_zipi8.t_state_1\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__18964\,
            I => \processor_zipi8.t_state_1\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__18961\,
            I => \processor_zipi8.t_state_1\
        );

    \I__3247\ : Odrv12
    port map (
            O => \N__18956\,
            I => \processor_zipi8.t_state_1\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__18953\,
            I => \processor_zipi8.t_state_1\
        );

    \I__3245\ : Odrv12
    port map (
            O => \N__18950\,
            I => \processor_zipi8.t_state_1\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__18935\,
            I => \processor_zipi8.decode4_strobes_enables_i.register_enable_type_0_cascade_\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__18932\,
            I => \N__18922\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__18931\,
            I => \N__18918\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__18930\,
            I => \N__18915\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__18929\,
            I => \N__18909\
        );

    \I__3239\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18903\
        );

    \I__3238\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18903\
        );

    \I__3237\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18898\
        );

    \I__3236\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18898\
        );

    \I__3235\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18895\
        );

    \I__3234\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18890\
        );

    \I__3233\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18890\
        );

    \I__3232\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18885\
        );

    \I__3231\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18885\
        );

    \I__3230\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18880\
        );

    \I__3229\ : InMux
    port map (
            O => \N__18912\,
            I => \N__18875\
        );

    \I__3228\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18875\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__18908\,
            I => \N__18871\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__18903\,
            I => \N__18868\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18863\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__18895\,
            I => \N__18863\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18858\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__18885\,
            I => \N__18858\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__18884\,
            I => \N__18855\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__18883\,
            I => \N__18852\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18849\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__18875\,
            I => \N__18846\
        );

    \I__3217\ : InMux
    port map (
            O => \N__18874\,
            I => \N__18841\
        );

    \I__3216\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18841\
        );

    \I__3215\ : Span4Mux_v
    port map (
            O => \N__18868\,
            I => \N__18836\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__18863\,
            I => \N__18836\
        );

    \I__3213\ : Span4Mux_s3_v
    port map (
            O => \N__18858\,
            I => \N__18833\
        );

    \I__3212\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18828\
        );

    \I__3211\ : InMux
    port map (
            O => \N__18852\,
            I => \N__18828\
        );

    \I__3210\ : Span4Mux_s2_h
    port map (
            O => \N__18849\,
            I => \N__18821\
        );

    \I__3209\ : Span4Mux_h
    port map (
            O => \N__18846\,
            I => \N__18821\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__18841\,
            I => \N__18821\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__18836\,
            I => instruction_17
        );

    \I__3206\ : Odrv4
    port map (
            O => \N__18833\,
            I => instruction_17
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__18828\,
            I => instruction_17
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__18821\,
            I => instruction_17
        );

    \I__3203\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18806\
        );

    \I__3202\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18806\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18806\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_22_3\
        );

    \I__3200\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18798\
        );

    \I__3199\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18794\
        );

    \I__3198\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18791\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__18798\,
            I => \N__18788\
        );

    \I__3196\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18785\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__18794\,
            I => \N__18778\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__18791\,
            I => \N__18778\
        );

    \I__3193\ : Span4Mux_v
    port map (
            O => \N__18788\,
            I => \N__18773\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18773\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__18784\,
            I => \N__18770\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__18783\,
            I => \N__18767\
        );

    \I__3189\ : Span4Mux_h
    port map (
            O => \N__18778\,
            I => \N__18762\
        );

    \I__3188\ : Span4Mux_h
    port map (
            O => \N__18773\,
            I => \N__18759\
        );

    \I__3187\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18750\
        );

    \I__3186\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18750\
        );

    \I__3185\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18750\
        );

    \I__3184\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18750\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__18762\,
            I => \processor_zipi8.sx_5\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__18759\,
            I => \processor_zipi8.sx_5\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__18750\,
            I => \processor_zipi8.sx_5\
        );

    \I__3180\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__18740\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_4\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__18737\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_4_cascade_\
        );

    \I__3177\ : InMux
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__18731\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_4\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__18728\,
            I => \N__18725\
        );

    \I__3174\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18719\
        );

    \I__3173\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18719\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__18719\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_4\
        );

    \I__3171\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18710\
        );

    \I__3170\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18710\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__18704\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_4\
        );

    \I__3166\ : InMux
    port map (
            O => \N__18701\,
            I => \N__18695\
        );

    \I__3165\ : InMux
    port map (
            O => \N__18700\,
            I => \N__18695\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__18689\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_4\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__18686\,
            I => \N__18682\
        );

    \I__3160\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18679\
        );

    \I__3159\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18676\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__18679\,
            I => \N__18671\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__18676\,
            I => \N__18671\
        );

    \I__3156\ : Span12Mux_s9_v
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__3155\ : Odrv12
    port map (
            O => \N__18668\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_4\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__18665\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_4_cascade_\
        );

    \I__3153\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__18659\,
            I => \N__18656\
        );

    \I__3151\ : Span4Mux_v
    port map (
            O => \N__18656\,
            I => \N__18653\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__18653\,
            I => \processor_zipi8.shift_rotate_result_4\
        );

    \I__3149\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__18641\,
            I => \processor_zipi8.spm_data_4\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__18638\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267_cascade_\
        );

    \I__3144\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18631\
        );

    \I__3143\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18628\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__18631\,
            I => \N__18623\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__18628\,
            I => \N__18623\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__18623\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_4\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__3138\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__18614\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_4\
        );

    \I__3136\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18607\
        );

    \I__3135\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18604\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__18607\,
            I => \N__18601\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__18604\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__18601\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4\
        );

    \I__3131\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__3128\ : Odrv4
    port map (
            O => \N__18587\,
            I => \processor_zipi8.shift_rotate_result_1\
        );

    \I__3127\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__18581\,
            I => \N__18578\
        );

    \I__3125\ : Span4Mux_h
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__18575\,
            I => \processor_zipi8.spm_data_1\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__18572\,
            I => \N__18568\
        );

    \I__3122\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18563\
        );

    \I__3121\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18563\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__3119\ : Odrv12
    port map (
            O => \N__18560\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_2\
        );

    \I__3118\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18553\
        );

    \I__3117\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18550\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18545\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18545\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__18542\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_2\
        );

    \I__3112\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__18536\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_2\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_2_cascade_\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__18530\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_2_cascade_\
        );

    \I__3108\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__18524\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_2\
        );

    \I__3106\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18517\
        );

    \I__3105\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18514\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__18517\,
            I => \N__18511\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__18514\,
            I => \N__18508\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__18511\,
            I => \N__18503\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__18508\,
            I => \N__18503\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__18500\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_3\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__3097\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__3095\ : Odrv12
    port map (
            O => \N__18488\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_am_1_3\
        );

    \I__3094\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18481\
        );

    \I__3093\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18478\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__18481\,
            I => \N__18475\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__18478\,
            I => \N__18472\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__18475\,
            I => \N__18469\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__18472\,
            I => \N__18466\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__18469\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__18466\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3\
        );

    \I__3086\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__18458\,
            I => \N__18454\
        );

    \I__3084\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18451\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__18454\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__18451\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2\
        );

    \I__3081\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18442\
        );

    \I__3080\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18439\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__18442\,
            I => \N__18436\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__18439\,
            I => \N__18433\
        );

    \I__3077\ : Span4Mux_h
    port map (
            O => \N__18436\,
            I => \N__18428\
        );

    \I__3076\ : Span4Mux_v
    port map (
            O => \N__18433\,
            I => \N__18428\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__18428\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_2\
        );

    \I__3074\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__18422\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_2\
        );

    \I__3072\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18413\
        );

    \I__3071\ : InMux
    port map (
            O => \N__18418\,
            I => \N__18413\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__18413\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_4\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__18410\,
            I => \N__18406\
        );

    \I__3068\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18401\
        );

    \I__3067\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18401\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__3065\ : Span4Mux_v
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__18395\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_4\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__18392\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_4_cascade_\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__18389\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_2_cascade_\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__3060\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18379\
        );

    \I__3059\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18376\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__18379\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__18376\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2\
        );

    \I__3056\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18365\
        );

    \I__3055\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18365\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__3053\ : Odrv4
    port map (
            O => \N__18362\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_2\
        );

    \I__3052\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__18356\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_bm_1_3\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__3049\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18344\
        );

    \I__3048\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18344\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__18344\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_3\
        );

    \I__3046\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18335\
        );

    \I__3045\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18335\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__3043\ : Odrv12
    port map (
            O => \N__18332\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_3\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__3041\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18322\
        );

    \I__3040\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18319\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__18322\,
            I => \N__18314\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__18319\,
            I => \N__18314\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__18311\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_5\
        );

    \I__3035\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18302\
        );

    \I__3034\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18302\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__18302\,
            I => \N__18299\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__18299\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_5\
        );

    \I__3031\ : InMux
    port map (
            O => \N__18296\,
            I => \N__18292\
        );

    \I__3030\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18289\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__18292\,
            I => \N__18286\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__18289\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5\
        );

    \I__3027\ : Odrv12
    port map (
            O => \N__18286\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_5_cascade_\
        );

    \I__3025\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__18275\,
            I => \N__18271\
        );

    \I__3023\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__3022\ : Odrv12
    port map (
            O => \N__18271\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__18268\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__18263\,
            I => \N__18260\
        );

    \I__3019\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__3017\ : Span4Mux_v
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__3016\ : Span4Mux_h
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__18248\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_179\
        );

    \I__3014\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18239\
        );

    \I__3013\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18239\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__18239\,
            I => \N__18236\
        );

    \I__3011\ : Span4Mux_v
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__18233\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_2\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__3008\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18223\
        );

    \I__3007\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18220\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__18223\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__18220\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__18215\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_2_cascade_\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__18212\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_3_cascade_\
        );

    \I__3002\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18205\
        );

    \I__3001\ : InMux
    port map (
            O => \N__18208\,
            I => \N__18202\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__18205\,
            I => \N__18199\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__18202\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__18199\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3\
        );

    \I__2997\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18188\
        );

    \I__2996\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18188\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__18185\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_3\
        );

    \I__2993\ : InMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__18179\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_3\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__18176\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_3_cascade_\
        );

    \I__2990\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18167\
        );

    \I__2989\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18167\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__18164\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_3\
        );

    \I__2986\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18155\
        );

    \I__2985\ : InMux
    port map (
            O => \N__18160\,
            I => \N__18155\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__18149\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_3\
        );

    \I__2981\ : InMux
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__18143\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_3\
        );

    \I__2979\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18136\
        );

    \I__2978\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__18136\,
            I => \N__18130\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__18133\,
            I => \N__18127\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__18130\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__18127\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__18122\,
            I => \N__18118\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__18121\,
            I => \N__18115\
        );

    \I__2971\ : InMux
    port map (
            O => \N__18118\,
            I => \N__18112\
        );

    \I__2970\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18109\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__18112\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__18109\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0\
        );

    \I__2967\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__2965\ : Span4Mux_s2_h
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__18092\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_5\
        );

    \I__2962\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__18086\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_3\
        );

    \I__2960\ : CEMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__2958\ : Span4Mux_v
    port map (
            O => \N__18077\,
            I => \N__18073\
        );

    \I__2957\ : CEMux
    port map (
            O => \N__18076\,
            I => \N__18070\
        );

    \I__2956\ : Span4Mux_h
    port map (
            O => \N__18073\,
            I => \N__18067\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__18070\,
            I => \N__18064\
        );

    \I__2954\ : Sp12to4
    port map (
            O => \N__18067\,
            I => \N__18059\
        );

    \I__2953\ : Span12Mux_s3_v
    port map (
            O => \N__18064\,
            I => \N__18059\
        );

    \I__2952\ : Odrv12
    port map (
            O => \N__18059\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe12\
        );

    \I__2951\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__18053\,
            I => \processor_zipi8.flags_i.use_zero_flagZ0\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \processor_zipi8.alu_result_0_cascade_\
        );

    \I__2948\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__18044\,
            I => \N__18039\
        );

    \I__2946\ : InMux
    port map (
            O => \N__18043\,
            I => \N__18034\
        );

    \I__2945\ : InMux
    port map (
            O => \N__18042\,
            I => \N__18034\
        );

    \I__2944\ : Span4Mux_v
    port map (
            O => \N__18039\,
            I => \N__18030\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__18034\,
            I => \N__18026\
        );

    \I__2942\ : InMux
    port map (
            O => \N__18033\,
            I => \N__18020\
        );

    \I__2941\ : Span4Mux_v
    port map (
            O => \N__18030\,
            I => \N__18017\
        );

    \I__2940\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18014\
        );

    \I__2939\ : Span4Mux_s2_v
    port map (
            O => \N__18026\,
            I => \N__18011\
        );

    \I__2938\ : InMux
    port map (
            O => \N__18025\,
            I => \N__18004\
        );

    \I__2937\ : InMux
    port map (
            O => \N__18024\,
            I => \N__18004\
        );

    \I__2936\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18004\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__18020\,
            I => \processor_zipi8.zero_flag\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__18017\,
            I => \processor_zipi8.zero_flag\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__18014\,
            I => \processor_zipi8.zero_flag\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__18011\,
            I => \processor_zipi8.zero_flag\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__18004\,
            I => \processor_zipi8.zero_flag\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__17993\,
            I => \N__17985\
        );

    \I__2929\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17981\
        );

    \I__2928\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17978\
        );

    \I__2927\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17975\
        );

    \I__2926\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17971\
        );

    \I__2925\ : InMux
    port map (
            O => \N__17988\,
            I => \N__17964\
        );

    \I__2924\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17964\
        );

    \I__2923\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17964\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__17981\,
            I => \N__17961\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__17978\,
            I => \N__17954\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__17975\,
            I => \N__17954\
        );

    \I__2919\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17951\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__17971\,
            I => \N__17946\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__17964\,
            I => \N__17946\
        );

    \I__2916\ : Span4Mux_h
    port map (
            O => \N__17961\,
            I => \N__17943\
        );

    \I__2915\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17938\
        );

    \I__2914\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17938\
        );

    \I__2913\ : Span4Mux_v
    port map (
            O => \N__17954\,
            I => \N__17931\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__17951\,
            I => \N__17931\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__17946\,
            I => \N__17931\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__17943\,
            I => \processor_zipi8.carry_flag\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__17938\,
            I => \processor_zipi8.carry_flag\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__17931\,
            I => \processor_zipi8.carry_flag\
        );

    \I__2907\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__17921\,
            I => \processor_zipi8.N_11_0\
        );

    \I__2905\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__17915\,
            I => \processor_zipi8.alu_result_1\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__17912\,
            I => \processor_zipi8.alu_result_2_cascade_\
        );

    \I__2902\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__17906\,
            I => \processor_zipi8.flags_i.zero_flag_3_0_0\
        );

    \I__2900\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17900\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__2898\ : Span4Mux_h
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__17894\,
            I => \processor_zipi8.flags_i.zero_flag_3_0_6\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__17891\,
            I => \N__17887\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__17890\,
            I => \N__17883\
        );

    \I__2894\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17872\
        );

    \I__2893\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17872\
        );

    \I__2892\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17872\
        );

    \I__2891\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17872\
        );

    \I__2890\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17868\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__17872\,
            I => \N__17865\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__17871\,
            I => \N__17862\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__17868\,
            I => \N__17854\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__17865\,
            I => \N__17851\
        );

    \I__2885\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17846\
        );

    \I__2884\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17841\
        );

    \I__2883\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17841\
        );

    \I__2882\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17834\
        );

    \I__2881\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17834\
        );

    \I__2880\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17834\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__17854\,
            I => \N__17831\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__17851\,
            I => \N__17828\
        );

    \I__2877\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17825\
        );

    \I__2876\ : InMux
    port map (
            O => \N__17849\,
            I => \N__17822\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__17846\,
            I => \N__17815\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17815\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__17834\,
            I => \N__17815\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__17831\,
            I => \processor_zipi8.pc_mode_2\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__17828\,
            I => \processor_zipi8.pc_mode_2\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__17825\,
            I => \processor_zipi8.pc_mode_2\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__17822\,
            I => \processor_zipi8.pc_mode_2\
        );

    \I__2868\ : Odrv12
    port map (
            O => \N__17815\,
            I => \processor_zipi8.pc_mode_2\
        );

    \I__2867\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17795\
        );

    \I__2866\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17786\
        );

    \I__2865\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17786\
        );

    \I__2864\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17786\
        );

    \I__2863\ : InMux
    port map (
            O => \N__17800\,
            I => \N__17786\
        );

    \I__2862\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17783\
        );

    \I__2861\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17780\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17777\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__17786\,
            I => \N__17768\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__17783\,
            I => \N__17763\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__17780\,
            I => \N__17763\
        );

    \I__2856\ : Span4Mux_v
    port map (
            O => \N__17777\,
            I => \N__17760\
        );

    \I__2855\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17755\
        );

    \I__2854\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17755\
        );

    \I__2853\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17746\
        );

    \I__2852\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17746\
        );

    \I__2851\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17746\
        );

    \I__2850\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17746\
        );

    \I__2849\ : Span4Mux_s1_h
    port map (
            O => \N__17768\,
            I => \N__17739\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__17763\,
            I => \N__17739\
        );

    \I__2847\ : Span4Mux_h
    port map (
            O => \N__17760\,
            I => \N__17739\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__17755\,
            I => \processor_zipi8.pc_mode_1\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__17746\,
            I => \processor_zipi8.pc_mode_1\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__17739\,
            I => \processor_zipi8.pc_mode_1\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__17732\,
            I => \N__17728\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__17731\,
            I => \N__17725\
        );

    \I__2841\ : CascadeBuf
    port map (
            O => \N__17728\,
            I => \N__17722\
        );

    \I__2840\ : CascadeBuf
    port map (
            O => \N__17725\,
            I => \N__17719\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__17722\,
            I => \N__17716\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__17719\,
            I => \N__17713\
        );

    \I__2837\ : CascadeBuf
    port map (
            O => \N__17716\,
            I => \N__17710\
        );

    \I__2836\ : CascadeBuf
    port map (
            O => \N__17713\,
            I => \N__17707\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__17710\,
            I => \N__17704\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__17707\,
            I => \N__17701\
        );

    \I__2833\ : CascadeBuf
    port map (
            O => \N__17704\,
            I => \N__17698\
        );

    \I__2832\ : CascadeBuf
    port map (
            O => \N__17701\,
            I => \N__17695\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__17698\,
            I => \N__17692\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__17695\,
            I => \N__17689\
        );

    \I__2829\ : CascadeBuf
    port map (
            O => \N__17692\,
            I => \N__17686\
        );

    \I__2828\ : CascadeBuf
    port map (
            O => \N__17689\,
            I => \N__17683\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__17686\,
            I => \N__17680\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__17683\,
            I => \N__17677\
        );

    \I__2825\ : CascadeBuf
    port map (
            O => \N__17680\,
            I => \N__17674\
        );

    \I__2824\ : CascadeBuf
    port map (
            O => \N__17677\,
            I => \N__17671\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__17674\,
            I => \N__17668\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__17671\,
            I => \N__17665\
        );

    \I__2821\ : CascadeBuf
    port map (
            O => \N__17668\,
            I => \N__17662\
        );

    \I__2820\ : CascadeBuf
    port map (
            O => \N__17665\,
            I => \N__17659\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__17662\,
            I => \N__17656\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__17659\,
            I => \N__17653\
        );

    \I__2817\ : CascadeBuf
    port map (
            O => \N__17656\,
            I => \N__17650\
        );

    \I__2816\ : CascadeBuf
    port map (
            O => \N__17653\,
            I => \N__17647\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__17650\,
            I => \N__17644\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__17647\,
            I => \N__17641\
        );

    \I__2813\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17636\
        );

    \I__2812\ : InMux
    port map (
            O => \N__17641\,
            I => \N__17633\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__17640\,
            I => \N__17630\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__17639\,
            I => \N__17627\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__17636\,
            I => \N__17624\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__17633\,
            I => \N__17621\
        );

    \I__2807\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17617\
        );

    \I__2806\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17614\
        );

    \I__2805\ : Span4Mux_s2_v
    port map (
            O => \N__17624\,
            I => \N__17609\
        );

    \I__2804\ : Span4Mux_s2_v
    port map (
            O => \N__17621\,
            I => \N__17609\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__17620\,
            I => \N__17605\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17602\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__17614\,
            I => \N__17599\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__17609\,
            I => \N__17596\
        );

    \I__2799\ : InMux
    port map (
            O => \N__17608\,
            I => \N__17593\
        );

    \I__2798\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17590\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__17602\,
            I => \N__17585\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__17599\,
            I => \N__17585\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__17596\,
            I => \N__17582\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__17593\,
            I => address_3
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__17590\,
            I => address_3
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__17585\,
            I => address_3
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__17582\,
            I => address_3
        );

    \I__2790\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__17570\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_3\
        );

    \I__2788\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__17564\,
            I => \N__17560\
        );

    \I__2786\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17557\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__17560\,
            I => \processor_zipi8.arith_carry_in_0\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__17557\,
            I => \processor_zipi8.arith_carry_in_0\
        );

    \I__2783\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__17546\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0\
        );

    \I__2780\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17539\
        );

    \I__2779\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17536\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17531\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__17536\,
            I => \N__17531\
        );

    \I__2776\ : Span4Mux_v
    port map (
            O => \N__17531\,
            I => \N__17527\
        );

    \I__2775\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17524\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__17527\,
            I => \processor_zipi8.returni_type_o_2\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__17524\,
            I => \processor_zipi8.returni_type_o_2\
        );

    \I__2772\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__17516\,
            I => \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_3\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__17513\,
            I => \processor_zipi8.decode4_strobes_enables_i.un9_flag_enable_type_cascade_\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__17510\,
            I => \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_0_cascade_\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__17507\,
            I => \N__17503\
        );

    \I__2767\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17500\
        );

    \I__2766\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17497\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__17500\,
            I => \N__17494\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__17497\,
            I => \N__17491\
        );

    \I__2763\ : Span4Mux_s1_h
    port map (
            O => \N__17494\,
            I => \N__17488\
        );

    \I__2762\ : Odrv12
    port map (
            O => \N__17491\,
            I => \processor_zipi8.flag_enable\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__17488\,
            I => \processor_zipi8.flag_enable\
        );

    \I__2760\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17480\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__17480\,
            I => \processor_zipi8.decode4_strobes_enables_i.spm_enable_value_1\
        );

    \I__2758\ : CEMux
    port map (
            O => \N__17477\,
            I => \N__17474\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__17474\,
            I => \N__17471\
        );

    \I__2756\ : Span4Mux_v
    port map (
            O => \N__17471\,
            I => \N__17468\
        );

    \I__2755\ : IoSpan4Mux
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__2754\ : IoSpan4Mux
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__2753\ : Span4Mux_s0_h
    port map (
            O => \N__17462\,
            I => \N__17459\
        );

    \I__2752\ : Span4Mux_h
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__2751\ : Odrv4
    port map (
            O => \N__17456\,
            I => \processor_zipi8.spm_enable\
        );

    \I__2750\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__17447\,
            I => \processor_zipi8.flags_i.carry_flag_value_1_0\
        );

    \I__2747\ : SRMux
    port map (
            O => \N__17444\,
            I => \N__17438\
        );

    \I__2746\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17435\
        );

    \I__2745\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17430\
        );

    \I__2744\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17430\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__17438\,
            I => \N__17426\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__17435\,
            I => \N__17420\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__17430\,
            I => \N__17420\
        );

    \I__2740\ : SRMux
    port map (
            O => \N__17429\,
            I => \N__17417\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__17426\,
            I => \N__17409\
        );

    \I__2738\ : SRMux
    port map (
            O => \N__17425\,
            I => \N__17406\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__17420\,
            I => \N__17395\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__17417\,
            I => \N__17395\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__17416\,
            I => \N__17391\
        );

    \I__2734\ : SRMux
    port map (
            O => \N__17415\,
            I => \N__17387\
        );

    \I__2733\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17380\
        );

    \I__2732\ : InMux
    port map (
            O => \N__17413\,
            I => \N__17380\
        );

    \I__2731\ : InMux
    port map (
            O => \N__17412\,
            I => \N__17380\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__17409\,
            I => \N__17374\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__17406\,
            I => \N__17374\
        );

    \I__2728\ : InMux
    port map (
            O => \N__17405\,
            I => \N__17365\
        );

    \I__2727\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17365\
        );

    \I__2726\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17365\
        );

    \I__2725\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17365\
        );

    \I__2724\ : SRMux
    port map (
            O => \N__17401\,
            I => \N__17362\
        );

    \I__2723\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17359\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__17395\,
            I => \N__17356\
        );

    \I__2721\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17351\
        );

    \I__2720\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17351\
        );

    \I__2719\ : SRMux
    port map (
            O => \N__17390\,
            I => \N__17348\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__17387\,
            I => \N__17345\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__17380\,
            I => \N__17342\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__17379\,
            I => \N__17336\
        );

    \I__2715\ : Span4Mux_s2_h
    port map (
            O => \N__17374\,
            I => \N__17331\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__17365\,
            I => \N__17331\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__17362\,
            I => \N__17322\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17322\
        );

    \I__2711\ : Sp12to4
    port map (
            O => \N__17356\,
            I => \N__17322\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__17351\,
            I => \N__17322\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__17348\,
            I => \N__17315\
        );

    \I__2708\ : Span4Mux_v
    port map (
            O => \N__17345\,
            I => \N__17315\
        );

    \I__2707\ : Span4Mux_v
    port map (
            O => \N__17342\,
            I => \N__17315\
        );

    \I__2706\ : InMux
    port map (
            O => \N__17341\,
            I => \N__17308\
        );

    \I__2705\ : InMux
    port map (
            O => \N__17340\,
            I => \N__17308\
        );

    \I__2704\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17308\
        );

    \I__2703\ : InMux
    port map (
            O => \N__17336\,
            I => \N__17305\
        );

    \I__2702\ : Span4Mux_s3_v
    port map (
            O => \N__17331\,
            I => \N__17302\
        );

    \I__2701\ : Span12Mux_s6_v
    port map (
            O => \N__17322\,
            I => \N__17299\
        );

    \I__2700\ : Span4Mux_h
    port map (
            O => \N__17315\,
            I => \N__17296\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__17308\,
            I => \processor_zipi8.internal_reset\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__17305\,
            I => \processor_zipi8.internal_reset\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__17302\,
            I => \processor_zipi8.internal_reset\
        );

    \I__2696\ : Odrv12
    port map (
            O => \N__17299\,
            I => \processor_zipi8.internal_reset\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__17296\,
            I => \processor_zipi8.internal_reset\
        );

    \I__2694\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17282\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__17282\,
            I => \N__17278\
        );

    \I__2692\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17275\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__17278\,
            I => \N__17270\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__17275\,
            I => \N__17270\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__17264\,
            I => \processor_zipi8.flags_i.N_69\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__17261\,
            I => \N__17256\
        );

    \I__2685\ : InMux
    port map (
            O => \N__17260\,
            I => \N__17252\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__17259\,
            I => \N__17248\
        );

    \I__2683\ : InMux
    port map (
            O => \N__17256\,
            I => \N__17245\
        );

    \I__2682\ : InMux
    port map (
            O => \N__17255\,
            I => \N__17242\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__17252\,
            I => \N__17239\
        );

    \I__2680\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17234\
        );

    \I__2679\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17234\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17231\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__17242\,
            I => \N__17227\
        );

    \I__2676\ : Sp12to4
    port map (
            O => \N__17239\,
            I => \N__17222\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__17234\,
            I => \N__17222\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__17231\,
            I => \N__17219\
        );

    \I__2673\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17216\
        );

    \I__2672\ : Span12Mux_s11_v
    port map (
            O => \N__17227\,
            I => \N__17211\
        );

    \I__2671\ : Span12Mux_s4_v
    port map (
            O => \N__17222\,
            I => \N__17211\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__17219\,
            I => \processor_zipi8.stack_pointer_3\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__17216\,
            I => \processor_zipi8.stack_pointer_3\
        );

    \I__2668\ : Odrv12
    port map (
            O => \N__17211\,
            I => \processor_zipi8.stack_pointer_3\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__17204\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_3_cascade_\
        );

    \I__2666\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__17198\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_3\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__17195\,
            I => \processor_zipi8.port_id_3_cascade_\
        );

    \I__2663\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__17189\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_3\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__17186\,
            I => \N__17182\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__17185\,
            I => \N__17179\
        );

    \I__2659\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__2658\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__17173\,
            I => \N__17167\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__17170\,
            I => \N__17163\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__17167\,
            I => \N__17160\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__17166\,
            I => \N__17157\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__17163\,
            I => \N__17152\
        );

    \I__2651\ : Sp12to4
    port map (
            O => \N__17160\,
            I => \N__17149\
        );

    \I__2650\ : InMux
    port map (
            O => \N__17157\,
            I => \N__17142\
        );

    \I__2649\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17142\
        );

    \I__2648\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17142\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__17152\,
            I => \processor_zipi8.port_id_3\
        );

    \I__2646\ : Odrv12
    port map (
            O => \N__17149\,
            I => \processor_zipi8.port_id_3\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__17142\,
            I => \processor_zipi8.port_id_3\
        );

    \I__2644\ : InMux
    port map (
            O => \N__17135\,
            I => \N__17132\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__17132\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_3\
        );

    \I__2642\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17110\
        );

    \I__2641\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17110\
        );

    \I__2640\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17110\
        );

    \I__2639\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17110\
        );

    \I__2638\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17110\
        );

    \I__2637\ : InMux
    port map (
            O => \N__17124\,
            I => \N__17103\
        );

    \I__2636\ : InMux
    port map (
            O => \N__17123\,
            I => \N__17103\
        );

    \I__2635\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17103\
        );

    \I__2634\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17097\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__17110\,
            I => \N__17092\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__17103\,
            I => \N__17092\
        );

    \I__2631\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17089\
        );

    \I__2630\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17084\
        );

    \I__2629\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17084\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__17097\,
            I => \N__17077\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__17092\,
            I => \N__17077\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__17089\,
            I => \N__17077\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__17084\,
            I => \N__17074\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__17077\,
            I => \N__17071\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__17074\,
            I => \N__17068\
        );

    \I__2622\ : Sp12to4
    port map (
            O => \N__17071\,
            I => \N__17065\
        );

    \I__2621\ : Sp12to4
    port map (
            O => \N__17068\,
            I => \N__17062\
        );

    \I__2620\ : Span12Mux_s2_h
    port map (
            O => \N__17065\,
            I => \N__17057\
        );

    \I__2619\ : Span12Mux_v
    port map (
            O => \N__17062\,
            I => \N__17057\
        );

    \I__2618\ : Odrv12
    port map (
            O => \N__17057\,
            I => instruction_3
        );

    \I__2617\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__17051\,
            I => \processor_zipi8.pc_vector_3\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__2614\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__17042\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_0\
        );

    \I__2612\ : InMux
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__17036\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4Z0Z_0\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__17033\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_cascade_\
        );

    \I__2609\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17027\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__17027\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__17024\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0_cascade_\
        );

    \I__2606\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__2604\ : Span4Mux_h
    port map (
            O => \N__17015\,
            I => \N__17011\
        );

    \I__2603\ : InMux
    port map (
            O => \N__17014\,
            I => \N__17008\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__17011\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__17008\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1\
        );

    \I__2600\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16997\
        );

    \I__2599\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16994\
        );

    \I__2598\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16989\
        );

    \I__2597\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16989\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16984\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__16994\,
            I => \N__16984\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__16989\,
            I => \N__16981\
        );

    \I__2593\ : Span4Mux_v
    port map (
            O => \N__16984\,
            I => \N__16976\
        );

    \I__2592\ : Span4Mux_v
    port map (
            O => \N__16981\,
            I => \N__16976\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__16973\,
            I => \N__16970\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__2588\ : Odrv4
    port map (
            O => \N__16967\,
            I => instruction_0
        );

    \I__2587\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__16961\,
            I => \N__16958\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__16955\,
            I => \processor_zipi8.register_bank_control_i.un1_bank_value\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__16952\,
            I => \processor_zipi8.register_bank_control_i.bank_0_1_cascade_\
        );

    \I__2582\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16945\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16948\,
            I => \N__16942\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__2578\ : Odrv12
    port map (
            O => \N__16939\,
            I => \processor_zipi8.sy_4\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__16936\,
            I => \processor_zipi8.sy_4\
        );

    \I__2576\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__16928\,
            I => \N__16925\
        );

    \I__2574\ : Span4Mux_h
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__2573\ : Span4Mux_s2_h
    port map (
            O => \N__16922\,
            I => \N__16919\
        );

    \I__2572\ : Odrv4
    port map (
            O => \N__16919\,
            I => \processor_zipi8.stack_i.stack_bank\
        );

    \I__2571\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__16913\,
            I => \processor_zipi8.shadow_bank\
        );

    \I__2569\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__16907\,
            I => \N__16904\
        );

    \I__2567\ : Span4Mux_h
    port map (
            O => \N__16904\,
            I => \N__16900\
        );

    \I__2566\ : InMux
    port map (
            O => \N__16903\,
            I => \N__16897\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__16900\,
            I => \processor_zipi8.un16_alu_mux_sel_value\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__16897\,
            I => \processor_zipi8.un16_alu_mux_sel_value\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__16892\,
            I => \processor_zipi8.un4_arith_logical_sel_cascade_\
        );

    \I__2562\ : InMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__2560\ : Span4Mux_s2_h
    port map (
            O => \N__16883\,
            I => \N__16880\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__16880\,
            I => \N__16876\
        );

    \I__2558\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16873\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__16876\,
            I => \processor_zipi8.alu_mux_sel_value_1\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__16873\,
            I => \processor_zipi8.alu_mux_sel_value_1\
        );

    \I__2555\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__16862\,
            I => \N__16858\
        );

    \I__2552\ : InMux
    port map (
            O => \N__16861\,
            I => \N__16855\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__16858\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__16855\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__16850\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2_cascade_\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__16847\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_0_cascade_\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__16844\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_0_cascade_\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__16841\,
            I => \N__16837\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__16840\,
            I => \N__16834\
        );

    \I__2544\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16831\
        );

    \I__2543\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16828\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__16831\,
            I => \N__16825\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__16828\,
            I => \N__16816\
        );

    \I__2540\ : Span4Mux_s3_h
    port map (
            O => \N__16825\,
            I => \N__16816\
        );

    \I__2539\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16811\
        );

    \I__2538\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16811\
        );

    \I__2537\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16806\
        );

    \I__2536\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16806\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__16816\,
            I => \processor_zipi8.port_id_0\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__16811\,
            I => \processor_zipi8.port_id_0\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__16806\,
            I => \processor_zipi8.port_id_0\
        );

    \I__2532\ : InMux
    port map (
            O => \N__16799\,
            I => \N__16793\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16798\,
            I => \N__16793\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__2529\ : Span4Mux_h
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__16787\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_6\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__16784\,
            I => \processor_zipi8.flags_i.carry_flag_value_1_1_cascade_\
        );

    \I__2526\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__16778\,
            I => \processor_zipi8.flags_i.parity_4\
        );

    \I__2524\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__16772\,
            I => \processor_zipi8.flags_i.carry_flag_RNOZ0Z_1\
        );

    \I__2522\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16765\
        );

    \I__2521\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16762\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__16765\,
            I => \processor_zipi8.flags_i.arith_carryZ0\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__16762\,
            I => \processor_zipi8.flags_i.arith_carryZ0\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__16757\,
            I => \N__16753\
        );

    \I__2517\ : InMux
    port map (
            O => \N__16756\,
            I => \N__16748\
        );

    \I__2516\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16748\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__16748\,
            I => \N__16745\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__2513\ : Span4Mux_h
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__16739\,
            I => \processor_zipi8.flags_i.shift_carryZ0\
        );

    \I__2511\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16733\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__16733\,
            I => \processor_zipi8.flags_i.carry_flag_value_1_0_0\
        );

    \I__2509\ : InMux
    port map (
            O => \N__16730\,
            I => \N__16727\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__16727\,
            I => \N__16724\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__16724\,
            I => \N__16721\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__16721\,
            I => \processor_zipi8.decode4_pc_statck_i.N_22_0\
        );

    \I__2505\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__16715\,
            I => \processor_zipi8.register_bank_control_i.un17_regbank_type_1\
        );

    \I__2503\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__16709\,
            I => \processor_zipi8.flags_i.un17_carry_flag_value_0\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__2500\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16698\
        );

    \I__2499\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16695\
        );

    \I__2498\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16691\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__16698\,
            I => \N__16686\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__16695\,
            I => \N__16686\
        );

    \I__2495\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16680\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__16691\,
            I => \N__16674\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__16686\,
            I => \N__16674\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__16685\,
            I => \N__16671\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__16684\,
            I => \N__16668\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__16683\,
            I => \N__16664\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__16680\,
            I => \N__16661\
        );

    \I__2488\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16658\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__16674\,
            I => \N__16655\
        );

    \I__2486\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16648\
        );

    \I__2485\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16648\
        );

    \I__2484\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16648\
        );

    \I__2483\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16645\
        );

    \I__2482\ : Odrv12
    port map (
            O => \N__16661\,
            I => \processor_zipi8.sx_7\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__16658\,
            I => \processor_zipi8.sx_7\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__16655\,
            I => \processor_zipi8.sx_7\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__16648\,
            I => \processor_zipi8.sx_7\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__16645\,
            I => \processor_zipi8.sx_7\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__16634\,
            I => \N__16627\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__16633\,
            I => \N__16624\
        );

    \I__2475\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16620\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \N__16616\
        );

    \I__2473\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16610\
        );

    \I__2472\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16610\
        );

    \I__2471\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16605\
        );

    \I__2470\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16605\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__16620\,
            I => \N__16602\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__16619\,
            I => \N__16599\
        );

    \I__2467\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16594\
        );

    \I__2466\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16594\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__16610\,
            I => \N__16589\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__16605\,
            I => \N__16589\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__16602\,
            I => \N__16586\
        );

    \I__2462\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16583\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__16594\,
            I => \N__16578\
        );

    \I__2460\ : Span4Mux_h
    port map (
            O => \N__16589\,
            I => \N__16578\
        );

    \I__2459\ : Span4Mux_s2_h
    port map (
            O => \N__16586\,
            I => \N__16575\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__16583\,
            I => \N__16572\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__16578\,
            I => \N__16569\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__16575\,
            I => \processor_zipi8.sx_6\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__16572\,
            I => \processor_zipi8.sx_6\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__16569\,
            I => \processor_zipi8.sx_6\
        );

    \I__2453\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16559\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__16559\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__16556\,
            I => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6_cascade_\
        );

    \I__2450\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16547\
        );

    \I__2449\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16547\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__16547\,
            I => \N__16544\
        );

    \I__2447\ : Odrv12
    port map (
            O => \N__16544\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_7\
        );

    \I__2446\ : InMux
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__16538\,
            I => \N__16534\
        );

    \I__2444\ : InMux
    port map (
            O => \N__16537\,
            I => \N__16531\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__16534\,
            I => \N__16526\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__16531\,
            I => \N__16526\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__16526\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_7\
        );

    \I__2440\ : CEMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__16514\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe15\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__16511\,
            I => \N__16507\
        );

    \I__2435\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16502\
        );

    \I__2434\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16502\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__16499\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_0\
        );

    \I__2431\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16490\
        );

    \I__2430\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16490\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__2428\ : Odrv12
    port map (
            O => \N__16487\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_5\
        );

    \I__2427\ : InMux
    port map (
            O => \N__16484\,
            I => \N__16478\
        );

    \I__2426\ : InMux
    port map (
            O => \N__16483\,
            I => \N__16478\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__16475\,
            I => \N__16472\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__16472\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_6\
        );

    \I__2422\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16463\
        );

    \I__2421\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16463\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__2419\ : Span4Mux_v
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__16457\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_7\
        );

    \I__2417\ : CEMux
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__16448\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe9\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__16445\,
            I => \N__16442\
        );

    \I__2413\ : InMux
    port map (
            O => \N__16442\,
            I => \N__16436\
        );

    \I__2412\ : InMux
    port map (
            O => \N__16441\,
            I => \N__16436\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__16430\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_6\
        );

    \I__2408\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16423\
        );

    \I__2407\ : InMux
    port map (
            O => \N__16426\,
            I => \N__16420\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__16423\,
            I => \N__16415\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__16420\,
            I => \N__16415\
        );

    \I__2404\ : Span4Mux_h
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__16412\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_7\
        );

    \I__2402\ : CEMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__16403\,
            I => \N__16400\
        );

    \I__2399\ : Span4Mux_s1_v
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__16397\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe13\
        );

    \I__2397\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16388\
        );

    \I__2396\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16388\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__16382\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_6\
        );

    \I__2392\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16375\
        );

    \I__2391\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16372\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__16375\,
            I => \N__16369\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16366\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__16369\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6\
        );

    \I__2387\ : Odrv12
    port map (
            O => \N__16366\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6\
        );

    \I__2386\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16357\
        );

    \I__2385\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16354\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__16357\,
            I => \N__16349\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__16354\,
            I => \N__16349\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__16349\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_6\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__16346\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_6_cascade_\
        );

    \I__2380\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16340\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__16340\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIK4HN1_6\
        );

    \I__2378\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16334\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__16331\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNII1NP1_6\
        );

    \I__2375\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16325\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__16325\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_6\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__16322\,
            I => \N__16319\
        );

    \I__2372\ : InMux
    port map (
            O => \N__16319\,
            I => \N__16316\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__16316\,
            I => \N__16313\
        );

    \I__2370\ : Span4Mux_h
    port map (
            O => \N__16313\,
            I => \N__16310\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__16310\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIGUSR1_6\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__16307\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7B4G8_6_cascade_\
        );

    \I__2367\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16301\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__16301\,
            I => \processor_zipi8.decode4_pc_statck_i.un3_pc_modeZ0\
        );

    \I__2365\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16295\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__16295\,
            I => \processor_zipi8.N_17_0\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__16292\,
            I => \N__16284\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__16291\,
            I => \N__16281\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__16290\,
            I => \N__16272\
        );

    \I__2360\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16265\
        );

    \I__2359\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16265\
        );

    \I__2358\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16262\
        );

    \I__2357\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16259\
        );

    \I__2356\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16256\
        );

    \I__2355\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16253\
        );

    \I__2354\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16246\
        );

    \I__2353\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16246\
        );

    \I__2352\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16246\
        );

    \I__2351\ : InMux
    port map (
            O => \N__16276\,
            I => \N__16237\
        );

    \I__2350\ : InMux
    port map (
            O => \N__16275\,
            I => \N__16237\
        );

    \I__2349\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16237\
        );

    \I__2348\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16237\
        );

    \I__2347\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16234\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__16265\,
            I => \N__16213\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__16262\,
            I => \N__16210\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__16259\,
            I => \N__16207\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__16256\,
            I => \N__16204\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__16253\,
            I => \N__16201\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__16246\,
            I => \N__16198\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__16237\,
            I => \N__16195\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__16234\,
            I => \N__16192\
        );

    \I__2338\ : CEMux
    port map (
            O => \N__16233\,
            I => \N__16139\
        );

    \I__2337\ : CEMux
    port map (
            O => \N__16232\,
            I => \N__16139\
        );

    \I__2336\ : CEMux
    port map (
            O => \N__16231\,
            I => \N__16139\
        );

    \I__2335\ : CEMux
    port map (
            O => \N__16230\,
            I => \N__16139\
        );

    \I__2334\ : CEMux
    port map (
            O => \N__16229\,
            I => \N__16139\
        );

    \I__2333\ : CEMux
    port map (
            O => \N__16228\,
            I => \N__16139\
        );

    \I__2332\ : CEMux
    port map (
            O => \N__16227\,
            I => \N__16139\
        );

    \I__2331\ : CEMux
    port map (
            O => \N__16226\,
            I => \N__16139\
        );

    \I__2330\ : CEMux
    port map (
            O => \N__16225\,
            I => \N__16139\
        );

    \I__2329\ : CEMux
    port map (
            O => \N__16224\,
            I => \N__16139\
        );

    \I__2328\ : CEMux
    port map (
            O => \N__16223\,
            I => \N__16139\
        );

    \I__2327\ : CEMux
    port map (
            O => \N__16222\,
            I => \N__16139\
        );

    \I__2326\ : CEMux
    port map (
            O => \N__16221\,
            I => \N__16139\
        );

    \I__2325\ : CEMux
    port map (
            O => \N__16220\,
            I => \N__16139\
        );

    \I__2324\ : CEMux
    port map (
            O => \N__16219\,
            I => \N__16139\
        );

    \I__2323\ : CEMux
    port map (
            O => \N__16218\,
            I => \N__16139\
        );

    \I__2322\ : CEMux
    port map (
            O => \N__16217\,
            I => \N__16139\
        );

    \I__2321\ : CEMux
    port map (
            O => \N__16216\,
            I => \N__16139\
        );

    \I__2320\ : Glb2LocalMux
    port map (
            O => \N__16213\,
            I => \N__16139\
        );

    \I__2319\ : Glb2LocalMux
    port map (
            O => \N__16210\,
            I => \N__16139\
        );

    \I__2318\ : Glb2LocalMux
    port map (
            O => \N__16207\,
            I => \N__16139\
        );

    \I__2317\ : Glb2LocalMux
    port map (
            O => \N__16204\,
            I => \N__16139\
        );

    \I__2316\ : Glb2LocalMux
    port map (
            O => \N__16201\,
            I => \N__16139\
        );

    \I__2315\ : Glb2LocalMux
    port map (
            O => \N__16198\,
            I => \N__16139\
        );

    \I__2314\ : Glb2LocalMux
    port map (
            O => \N__16195\,
            I => \N__16139\
        );

    \I__2313\ : Glb2LocalMux
    port map (
            O => \N__16192\,
            I => \N__16139\
        );

    \I__2312\ : GlobalMux
    port map (
            O => \N__16139\,
            I => \N__16136\
        );

    \I__2311\ : gio2CtrlBuf
    port map (
            O => \N__16136\,
            I => bram_enable_g
        );

    \I__2310\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16130\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__16130\,
            I => \N__16127\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__16127\,
            I => \processor_zipi8.flags_i.m104Z0Z_2\
        );

    \I__2307\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16120\
        );

    \I__2306\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16117\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__16120\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__16117\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6\
        );

    \I__2303\ : InMux
    port map (
            O => \N__16112\,
            I => \N__16108\
        );

    \I__2302\ : InMux
    port map (
            O => \N__16111\,
            I => \N__16105\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__16108\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__16105\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__16100\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_6_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__16097\,
            I => \N__16094\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__16094\,
            I => \N__16090\
        );

    \I__2296\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16087\
        );

    \I__2295\ : Span4Mux_h
    port map (
            O => \N__16090\,
            I => \N__16082\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__16087\,
            I => \N__16082\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__16082\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_6\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__16079\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI44F42_6_cascade_\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__16076\,
            I => \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_1_cascade_\
        );

    \I__2290\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16070\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__16070\,
            I => \N__16067\
        );

    \I__2288\ : Odrv12
    port map (
            O => \N__16067\,
            I => \processor_zipi8.shift_rotate_result_2\
        );

    \I__2287\ : InMux
    port map (
            O => \N__16064\,
            I => \N__16061\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__2285\ : Span4Mux_v
    port map (
            O => \N__16058\,
            I => \N__16055\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__16055\,
            I => \processor_zipi8.spm_data_2\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__16052\,
            I => \processor_zipi8.register_bank_control_i.un31_regbank_type_3_cascade_\
        );

    \I__2282\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16046\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__2280\ : Odrv12
    port map (
            O => \N__16043\,
            I => \processor_zipi8.register_bank_control_i.un31_regbank_type\
        );

    \I__2279\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16037\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__16037\,
            I => \N__16034\
        );

    \I__2277\ : Odrv12
    port map (
            O => \N__16034\,
            I => \processor_zipi8.shift_rotate_result_0\
        );

    \I__2276\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16028\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__16025\,
            I => \N__16022\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__16019\,
            I => \processor_zipi8.spm_data_0\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__16016\,
            I => \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_0_cascade_\
        );

    \I__2270\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16007\
        );

    \I__2269\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16007\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__16001\,
            I => \processor_zipi8.pc_mode_2_0_0\
        );

    \I__2265\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__2263\ : Odrv12
    port map (
            O => \N__15992\,
            I => \processor_zipi8.pc_vector_2\
        );

    \I__2262\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__15983\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_2\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__2258\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15971\
        );

    \I__2257\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15971\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15967\
        );

    \I__2255\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15964\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__15967\,
            I => \processor_zipi8.program_counter_i.half_pc_0_2\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__15964\,
            I => \processor_zipi8.program_counter_i.half_pc_0_2\
        );

    \I__2252\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15949\
        );

    \I__2251\ : InMux
    port map (
            O => \N__15958\,
            I => \N__15949\
        );

    \I__2250\ : InMux
    port map (
            O => \N__15957\,
            I => \N__15946\
        );

    \I__2249\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15941\
        );

    \I__2248\ : InMux
    port map (
            O => \N__15955\,
            I => \N__15941\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__15954\,
            I => \N__15929\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15921\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__15946\,
            I => \N__15921\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__15941\,
            I => \N__15918\
        );

    \I__2243\ : InMux
    port map (
            O => \N__15940\,
            I => \N__15913\
        );

    \I__2242\ : InMux
    port map (
            O => \N__15939\,
            I => \N__15913\
        );

    \I__2241\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15910\
        );

    \I__2240\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15903\
        );

    \I__2239\ : InMux
    port map (
            O => \N__15936\,
            I => \N__15903\
        );

    \I__2238\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15903\
        );

    \I__2237\ : InMux
    port map (
            O => \N__15934\,
            I => \N__15888\
        );

    \I__2236\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15888\
        );

    \I__2235\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15888\
        );

    \I__2234\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15888\
        );

    \I__2233\ : InMux
    port map (
            O => \N__15928\,
            I => \N__15888\
        );

    \I__2232\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15888\
        );

    \I__2231\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15888\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__15921\,
            I => \N__15885\
        );

    \I__2229\ : Span4Mux_h
    port map (
            O => \N__15918\,
            I => \N__15882\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__15913\,
            I => \processor_zipi8.program_counter_i.un3_half_pcZ0\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__15910\,
            I => \processor_zipi8.program_counter_i.un3_half_pcZ0\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__15903\,
            I => \processor_zipi8.program_counter_i.un3_half_pcZ0\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__15888\,
            I => \processor_zipi8.program_counter_i.un3_half_pcZ0\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__15885\,
            I => \processor_zipi8.program_counter_i.un3_half_pcZ0\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__15882\,
            I => \processor_zipi8.program_counter_i.un3_half_pcZ0\
        );

    \I__2222\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15866\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15862\
        );

    \I__2220\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15859\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__15862\,
            I => \processor_zipi8.program_counter_i.half_pc_0_3\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__15859\,
            I => \processor_zipi8.program_counter_i.half_pc_0_3\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__15854\,
            I => \processor_zipi8.un16_alu_mux_sel_value_cascade_\
        );

    \I__2216\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15848\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__15848\,
            I => \processor_zipi8.decode4_strobes_enables_i.un23_flag_enable_type\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__15845\,
            I => \processor_zipi8.pc_vector_0_cascade_\
        );

    \I__2213\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15836\
        );

    \I__2212\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15836\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__15836\,
            I => \N__15833\
        );

    \I__2210\ : Span4Mux_h
    port map (
            O => \N__15833\,
            I => \N__15830\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__15830\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_0\
        );

    \I__2208\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15823\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__15826\,
            I => \N__15820\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__15823\,
            I => \N__15817\
        );

    \I__2205\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15814\
        );

    \I__2204\ : Span4Mux_s3_h
    port map (
            O => \N__15817\,
            I => \N__15811\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__15814\,
            I => \N__15808\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__15811\,
            I => \processor_zipi8.flags_i.i14_mux\
        );

    \I__2201\ : Odrv12
    port map (
            O => \N__15808\,
            I => \processor_zipi8.flags_i.i14_mux\
        );

    \I__2200\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15799\
        );

    \I__2199\ : InMux
    port map (
            O => \N__15802\,
            I => \N__15796\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__15799\,
            I => \N__15793\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__15796\,
            I => \N__15790\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__15793\,
            I => \N__15787\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__15790\,
            I => \N__15784\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__15787\,
            I => \processor_zipi8.flags_i.i14_mux_0\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__15784\,
            I => \processor_zipi8.flags_i.i14_mux_0\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__2191\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__15770\,
            I => \processor_zipi8.zero_flag_RNIC4FP9\
        );

    \I__2188\ : CEMux
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__15764\,
            I => \N__15759\
        );

    \I__2186\ : CEMux
    port map (
            O => \N__15763\,
            I => \N__15755\
        );

    \I__2185\ : CEMux
    port map (
            O => \N__15762\,
            I => \N__15752\
        );

    \I__2184\ : Span4Mux_v
    port map (
            O => \N__15759\,
            I => \N__15749\
        );

    \I__2183\ : CEMux
    port map (
            O => \N__15758\,
            I => \N__15746\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__15755\,
            I => \N__15743\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__15752\,
            I => \N__15740\
        );

    \I__2180\ : Span4Mux_s1_h
    port map (
            O => \N__15749\,
            I => \N__15737\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15734\
        );

    \I__2178\ : Span4Mux_s2_h
    port map (
            O => \N__15743\,
            I => \N__15729\
        );

    \I__2177\ : Span4Mux_s2_h
    port map (
            O => \N__15740\,
            I => \N__15729\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__15737\,
            I => \processor_zipi8.program_counter_i.t_state_0_1\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__15734\,
            I => \processor_zipi8.program_counter_i.t_state_0_1\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__15729\,
            I => \processor_zipi8.program_counter_i.t_state_0_1\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__15722\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_1_cascade_\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__15719\,
            I => \processor_zipi8.program_counter_i.half_pc_0_1_cascade_\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__15716\,
            I => \N__15712\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \N__15709\
        );

    \I__2169\ : CascadeBuf
    port map (
            O => \N__15712\,
            I => \N__15706\
        );

    \I__2168\ : CascadeBuf
    port map (
            O => \N__15709\,
            I => \N__15703\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__15706\,
            I => \N__15700\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__15703\,
            I => \N__15697\
        );

    \I__2165\ : CascadeBuf
    port map (
            O => \N__15700\,
            I => \N__15694\
        );

    \I__2164\ : CascadeBuf
    port map (
            O => \N__15697\,
            I => \N__15691\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__15694\,
            I => \N__15688\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__15691\,
            I => \N__15685\
        );

    \I__2161\ : CascadeBuf
    port map (
            O => \N__15688\,
            I => \N__15682\
        );

    \I__2160\ : CascadeBuf
    port map (
            O => \N__15685\,
            I => \N__15679\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__15682\,
            I => \N__15676\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__15679\,
            I => \N__15673\
        );

    \I__2157\ : CascadeBuf
    port map (
            O => \N__15676\,
            I => \N__15670\
        );

    \I__2156\ : CascadeBuf
    port map (
            O => \N__15673\,
            I => \N__15667\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__15670\,
            I => \N__15664\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__15667\,
            I => \N__15661\
        );

    \I__2153\ : CascadeBuf
    port map (
            O => \N__15664\,
            I => \N__15658\
        );

    \I__2152\ : CascadeBuf
    port map (
            O => \N__15661\,
            I => \N__15655\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__15658\,
            I => \N__15652\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__15655\,
            I => \N__15649\
        );

    \I__2149\ : CascadeBuf
    port map (
            O => \N__15652\,
            I => \N__15646\
        );

    \I__2148\ : CascadeBuf
    port map (
            O => \N__15649\,
            I => \N__15643\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__15646\,
            I => \N__15640\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__15643\,
            I => \N__15637\
        );

    \I__2145\ : CascadeBuf
    port map (
            O => \N__15640\,
            I => \N__15634\
        );

    \I__2144\ : CascadeBuf
    port map (
            O => \N__15637\,
            I => \N__15631\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__15634\,
            I => \N__15627\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__15631\,
            I => \N__15624\
        );

    \I__2141\ : InMux
    port map (
            O => \N__15630\,
            I => \N__15621\
        );

    \I__2140\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15618\
        );

    \I__2139\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15615\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__15621\,
            I => \N__15612\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__15618\,
            I => \N__15606\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__15615\,
            I => \N__15603\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__15612\,
            I => \N__15599\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__15611\,
            I => \N__15596\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__15610\,
            I => \N__15593\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__15609\,
            I => \N__15590\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__15606\,
            I => \N__15587\
        );

    \I__2130\ : Span4Mux_s3_h
    port map (
            O => \N__15603\,
            I => \N__15584\
        );

    \I__2129\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15581\
        );

    \I__2128\ : Sp12to4
    port map (
            O => \N__15599\,
            I => \N__15578\
        );

    \I__2127\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15575\
        );

    \I__2126\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15572\
        );

    \I__2125\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15569\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__15587\,
            I => \N__15566\
        );

    \I__2123\ : Span4Mux_h
    port map (
            O => \N__15584\,
            I => \N__15563\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__15581\,
            I => address_1
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__15578\,
            I => address_1
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__15575\,
            I => address_1
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__15572\,
            I => address_1
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__15569\,
            I => address_1
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__15566\,
            I => address_1
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__15563\,
            I => address_1
        );

    \I__2115\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15545\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__15545\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__15542\,
            I => \N__15538\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__15541\,
            I => \N__15535\
        );

    \I__2111\ : CascadeBuf
    port map (
            O => \N__15538\,
            I => \N__15532\
        );

    \I__2110\ : CascadeBuf
    port map (
            O => \N__15535\,
            I => \N__15529\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__15532\,
            I => \N__15526\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__15529\,
            I => \N__15523\
        );

    \I__2107\ : CascadeBuf
    port map (
            O => \N__15526\,
            I => \N__15520\
        );

    \I__2106\ : CascadeBuf
    port map (
            O => \N__15523\,
            I => \N__15517\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__15520\,
            I => \N__15514\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__15517\,
            I => \N__15511\
        );

    \I__2103\ : CascadeBuf
    port map (
            O => \N__15514\,
            I => \N__15508\
        );

    \I__2102\ : CascadeBuf
    port map (
            O => \N__15511\,
            I => \N__15505\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__15508\,
            I => \N__15502\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__15505\,
            I => \N__15499\
        );

    \I__2099\ : CascadeBuf
    port map (
            O => \N__15502\,
            I => \N__15496\
        );

    \I__2098\ : CascadeBuf
    port map (
            O => \N__15499\,
            I => \N__15493\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__15496\,
            I => \N__15490\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__15493\,
            I => \N__15487\
        );

    \I__2095\ : CascadeBuf
    port map (
            O => \N__15490\,
            I => \N__15484\
        );

    \I__2094\ : CascadeBuf
    port map (
            O => \N__15487\,
            I => \N__15481\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__15484\,
            I => \N__15478\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__15481\,
            I => \N__15475\
        );

    \I__2091\ : CascadeBuf
    port map (
            O => \N__15478\,
            I => \N__15472\
        );

    \I__2090\ : CascadeBuf
    port map (
            O => \N__15475\,
            I => \N__15469\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__15472\,
            I => \N__15466\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__15469\,
            I => \N__15463\
        );

    \I__2087\ : CascadeBuf
    port map (
            O => \N__15466\,
            I => \N__15460\
        );

    \I__2086\ : CascadeBuf
    port map (
            O => \N__15463\,
            I => \N__15457\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__15460\,
            I => \N__15454\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__15457\,
            I => \N__15451\
        );

    \I__2083\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15445\
        );

    \I__2082\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15442\
        );

    \I__2081\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15438\
        );

    \I__2080\ : InMux
    port map (
            O => \N__15449\,
            I => \N__15434\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__15448\,
            I => \N__15431\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__15445\,
            I => \N__15426\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__15442\,
            I => \N__15426\
        );

    \I__2076\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15423\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__15438\,
            I => \N__15420\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__15437\,
            I => \N__15417\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__15434\,
            I => \N__15414\
        );

    \I__2072\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15411\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__15426\,
            I => \N__15408\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__15423\,
            I => \N__15403\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__15420\,
            I => \N__15403\
        );

    \I__2068\ : InMux
    port map (
            O => \N__15417\,
            I => \N__15400\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__15414\,
            I => \N__15393\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__15411\,
            I => \N__15393\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__15408\,
            I => \N__15393\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__15403\,
            I => address_0
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__15400\,
            I => address_0
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__15393\,
            I => address_0
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__15386\,
            I => \N__15383\
        );

    \I__2060\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15380\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__2058\ : Span4Mux_s3_h
    port map (
            O => \N__15377\,
            I => \N__15374\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__15374\,
            I => \processor_zipi8.zero_flag_RNIL8RB5\
        );

    \I__2056\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15364\
        );

    \I__2055\ : InMux
    port map (
            O => \N__15370\,
            I => \N__15364\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__15369\,
            I => \N__15361\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__15364\,
            I => \N__15358\
        );

    \I__2052\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15355\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__15358\,
            I => \processor_zipi8.program_counter_i.half_pc_0_1\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__15355\,
            I => \processor_zipi8.program_counter_i.half_pc_0_1\
        );

    \I__2049\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15342\
        );

    \I__2048\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15342\
        );

    \I__2047\ : InMux
    port map (
            O => \N__15348\,
            I => \N__15337\
        );

    \I__2046\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15337\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__15342\,
            I => \processor_zipi8.program_counter_i.carry_pc_4_0\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__15337\,
            I => \processor_zipi8.program_counter_i.carry_pc_4_0\
        );

    \I__2043\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15326\
        );

    \I__2042\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15326\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__15326\,
            I => \N__15323\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__15323\,
            I => \processor_zipi8.program_counter_i.carry_pc_22_3\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__2038\ : CascadeBuf
    port map (
            O => \N__15317\,
            I => \N__15314\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__15314\,
            I => \N__15310\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__15313\,
            I => \N__15307\
        );

    \I__2035\ : CascadeBuf
    port map (
            O => \N__15310\,
            I => \N__15304\
        );

    \I__2034\ : CascadeBuf
    port map (
            O => \N__15307\,
            I => \N__15301\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__15304\,
            I => \N__15298\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__15301\,
            I => \N__15295\
        );

    \I__2031\ : CascadeBuf
    port map (
            O => \N__15298\,
            I => \N__15292\
        );

    \I__2030\ : CascadeBuf
    port map (
            O => \N__15295\,
            I => \N__15289\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__15292\,
            I => \N__15286\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__15289\,
            I => \N__15283\
        );

    \I__2027\ : CascadeBuf
    port map (
            O => \N__15286\,
            I => \N__15280\
        );

    \I__2026\ : CascadeBuf
    port map (
            O => \N__15283\,
            I => \N__15277\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__15280\,
            I => \N__15274\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__15277\,
            I => \N__15271\
        );

    \I__2023\ : CascadeBuf
    port map (
            O => \N__15274\,
            I => \N__15268\
        );

    \I__2022\ : CascadeBuf
    port map (
            O => \N__15271\,
            I => \N__15265\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__15268\,
            I => \N__15262\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__15265\,
            I => \N__15259\
        );

    \I__2019\ : CascadeBuf
    port map (
            O => \N__15262\,
            I => \N__15256\
        );

    \I__2018\ : CascadeBuf
    port map (
            O => \N__15259\,
            I => \N__15253\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__15256\,
            I => \N__15250\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__15253\,
            I => \N__15247\
        );

    \I__2015\ : CascadeBuf
    port map (
            O => \N__15250\,
            I => \N__15244\
        );

    \I__2014\ : CascadeBuf
    port map (
            O => \N__15247\,
            I => \N__15241\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__15244\,
            I => \N__15238\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__15241\,
            I => \N__15235\
        );

    \I__2011\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15231\
        );

    \I__2010\ : CascadeBuf
    port map (
            O => \N__15235\,
            I => \N__15228\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__15234\,
            I => \N__15224\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__15231\,
            I => \N__15221\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__15228\,
            I => \N__15218\
        );

    \I__2006\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15215\
        );

    \I__2005\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15211\
        );

    \I__2004\ : Span4Mux_s1_v
    port map (
            O => \N__15221\,
            I => \N__15208\
        );

    \I__2003\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15205\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__15215\,
            I => \N__15201\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__15214\,
            I => \N__15198\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__15211\,
            I => \N__15195\
        );

    \I__1999\ : Sp12to4
    port map (
            O => \N__15208\,
            I => \N__15190\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__15205\,
            I => \N__15190\
        );

    \I__1997\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15187\
        );

    \I__1996\ : Span4Mux_s3_h
    port map (
            O => \N__15201\,
            I => \N__15184\
        );

    \I__1995\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15181\
        );

    \I__1994\ : Sp12to4
    port map (
            O => \N__15195\,
            I => \N__15176\
        );

    \I__1993\ : Span12Mux_s8_h
    port map (
            O => \N__15190\,
            I => \N__15176\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__15187\,
            I => address_2
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__15184\,
            I => address_2
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__15181\,
            I => address_2
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__15176\,
            I => address_2
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__15167\,
            I => \N__15162\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__15166\,
            I => \N__15159\
        );

    \I__1986\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15154\
        );

    \I__1985\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15151\
        );

    \I__1984\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15148\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__15158\,
            I => \N__15145\
        );

    \I__1982\ : InMux
    port map (
            O => \N__15157\,
            I => \N__15141\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__15154\,
            I => \N__15136\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__15151\,
            I => \N__15136\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__15148\,
            I => \N__15133\
        );

    \I__1978\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15128\
        );

    \I__1977\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15128\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__15141\,
            I => \N__15125\
        );

    \I__1975\ : Span4Mux_s2_v
    port map (
            O => \N__15136\,
            I => \N__15122\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__15133\,
            I => \processor_zipi8.stack_pointer_4\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__15128\,
            I => \processor_zipi8.stack_pointer_4\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__15125\,
            I => \processor_zipi8.stack_pointer_4\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__15122\,
            I => \processor_zipi8.stack_pointer_4\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__1969\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15106\
        );

    \I__1968\ : InMux
    port map (
            O => \N__15109\,
            I => \N__15103\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__15106\,
            I => \N__15097\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15097\
        );

    \I__1965\ : InMux
    port map (
            O => \N__15102\,
            I => \N__15094\
        );

    \I__1964\ : Span4Mux_h
    port map (
            O => \N__15097\,
            I => \N__15091\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__15094\,
            I => \N__15088\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__15091\,
            I => \processor_zipi8.flags_i.N_34\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__15088\,
            I => \processor_zipi8.flags_i.N_34\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__15083\,
            I => \processor_zipi8.port_id_0_cascade_\
        );

    \I__1959\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__15071\,
            I => \processor_zipi8.stack_memory_0\
        );

    \I__1955\ : InMux
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__15065\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_0\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__15062\,
            I => \N__15059\
        );

    \I__1952\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15056\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__15056\,
            I => \N__15053\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__15053\,
            I => \processor_zipi8.pc_vector_0\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__15050\,
            I => \N__15046\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__15049\,
            I => \N__15042\
        );

    \I__1947\ : InMux
    port map (
            O => \N__15046\,
            I => \N__15039\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__15045\,
            I => \N__15036\
        );

    \I__1945\ : InMux
    port map (
            O => \N__15042\,
            I => \N__15031\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__15039\,
            I => \N__15028\
        );

    \I__1943\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15025\
        );

    \I__1942\ : InMux
    port map (
            O => \N__15035\,
            I => \N__15020\
        );

    \I__1941\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15020\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__15031\,
            I => \processor_zipi8.port_id_2\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__15028\,
            I => \processor_zipi8.port_id_2\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__15025\,
            I => \processor_zipi8.port_id_2\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__15020\,
            I => \processor_zipi8.port_id_2\
        );

    \I__1936\ : InMux
    port map (
            O => \N__15011\,
            I => \N__15008\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__15008\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_2\
        );

    \I__1934\ : InMux
    port map (
            O => \N__15005\,
            I => \N__15002\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__15002\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_2\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__14999\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_2_cascade_\
        );

    \I__1931\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__14993\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_2\
        );

    \I__1929\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14987\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__1927\ : Span4Mux_h
    port map (
            O => \N__14984\,
            I => \N__14981\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__14981\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_2\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__14978\,
            I => \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_0_cascade_\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__14975\,
            I => \N__14970\
        );

    \I__1923\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14961\
        );

    \I__1922\ : InMux
    port map (
            O => \N__14973\,
            I => \N__14961\
        );

    \I__1921\ : InMux
    port map (
            O => \N__14970\,
            I => \N__14961\
        );

    \I__1920\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14958\
        );

    \I__1919\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14955\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__14961\,
            I => \N__14948\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__14958\,
            I => \N__14948\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__14955\,
            I => \N__14948\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__14948\,
            I => \N__14945\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__14945\,
            I => \N__14942\
        );

    \I__1913\ : Span4Mux_h
    port map (
            O => \N__14942\,
            I => \N__14939\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__14939\,
            I => instruction_2
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__14936\,
            I => \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_1_cascade_\
        );

    \I__1910\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14927\
        );

    \I__1909\ : InMux
    port map (
            O => \N__14932\,
            I => \N__14927\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__14924\,
            I => \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_0\
        );

    \I__1906\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14918\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__1904\ : Odrv12
    port map (
            O => \N__14915\,
            I => \processor_zipi8.shift_rotate_result_6\
        );

    \I__1903\ : InMux
    port map (
            O => \N__14912\,
            I => \N__14909\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__14909\,
            I => \N__14906\
        );

    \I__1901\ : Span4Mux_s3_h
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__14903\,
            I => \processor_zipi8.shift_rotate_result_5\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \processor_zipi8.port_id_2_cascade_\
        );

    \I__1898\ : CEMux
    port map (
            O => \N__14897\,
            I => \N__14894\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__1896\ : Span4Mux_s3_h
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__14888\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe11\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__14885\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212_cascade_\
        );

    \I__1893\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__14879\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_0\
        );

    \I__1891\ : CEMux
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__1889\ : Span4Mux_s3_h
    port map (
            O => \N__14870\,
            I => \N__14867\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__14867\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe8\
        );

    \I__1887\ : CEMux
    port map (
            O => \N__14864\,
            I => \N__14860\
        );

    \I__1886\ : CEMux
    port map (
            O => \N__14863\,
            I => \N__14857\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__14860\,
            I => \N__14854\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__14857\,
            I => \N__14851\
        );

    \I__1883\ : Span4Mux_s1_v
    port map (
            O => \N__14854\,
            I => \N__14848\
        );

    \I__1882\ : Span4Mux_s3_h
    port map (
            O => \N__14851\,
            I => \N__14845\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__14848\,
            I => \N__14842\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__14845\,
            I => \N__14839\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__14842\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__14839\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__14834\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268_cascade_\
        );

    \I__1876\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14828\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__14828\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_6\
        );

    \I__1874\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14819\
        );

    \I__1873\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14819\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__14819\,
            I => \N__14816\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__14813\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_0\
        );

    \I__1869\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14804\
        );

    \I__1868\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14804\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__1866\ : Span4Mux_h
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__14798\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_0\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__14795\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_0_cascade_\
        );

    \I__1863\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14786\
        );

    \I__1862\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14786\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__1860\ : Sp12to4
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__1859\ : Odrv12
    port map (
            O => \N__14780\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_0\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__14777\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_0_cascade_\
        );

    \I__1857\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__14771\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_0\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__14768\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_0_cascade_\
        );

    \I__1854\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14762\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__14762\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_0\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__14759\,
            I => \processor_zipi8.flags_i.m68_ns_1_cascade_\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__14756\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_6_cascade_\
        );

    \I__1850\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14750\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__14747\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_6\
        );

    \I__1847\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__14741\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_6\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__14738\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_6_cascade_\
        );

    \I__1844\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__14732\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_6\
        );

    \I__1842\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14723\
        );

    \I__1840\ : Span4Mux_h
    port map (
            O => \N__14723\,
            I => \N__14720\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__14720\,
            I => \processor_zipi8.spm_data_6\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__14717\,
            I => \processor_zipi8.flags_i.N_1235_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__14711\,
            I => \processor_zipi8.flags_i.zero_flag_RNI89VZ0Z91\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__1834\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14702\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__14702\,
            I => \processor_zipi8.flags_i.N_1239\
        );

    \I__1832\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14696\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__14696\,
            I => \processor_zipi8.flags_i.N_124_mux\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__14693\,
            I => \processor_zipi8.flags_i.N_1241_cascade_\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__14690\,
            I => \N__14687\
        );

    \I__1828\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__14678\,
            I => \processor_zipi8.zero_flag_RNIDS654\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__1823\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__1820\ : Span4Mux_v
    port map (
            O => \N__14663\,
            I => \N__14654\
        );

    \I__1819\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14651\
        );

    \I__1818\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14648\
        );

    \I__1817\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14643\
        );

    \I__1816\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14643\
        );

    \I__1815\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14640\
        );

    \I__1814\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14637\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__14654\,
            I => \processor_zipi8.stack_pointer_1\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__14651\,
            I => \processor_zipi8.stack_pointer_1\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__14648\,
            I => \processor_zipi8.stack_pointer_1\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__14643\,
            I => \processor_zipi8.stack_pointer_1\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__14640\,
            I => \processor_zipi8.stack_pointer_1\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__14637\,
            I => \processor_zipi8.stack_pointer_1\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__1806\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__14618\,
            I => \processor_zipi8.flags_i.m75_amZ0\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__14615\,
            I => \processor_zipi8.flags_i.m75_amZ0_cascade_\
        );

    \I__1803\ : InMux
    port map (
            O => \N__14612\,
            I => \N__14606\
        );

    \I__1802\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14606\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__14606\,
            I => \processor_zipi8.flags_i.zero_flag_RNI3VCZ0Z94\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__1799\ : InMux
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__14591\,
            I => \processor_zipi8.zero_flag_RNI5GK75\
        );

    \I__1795\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__14585\,
            I => \processor_zipi8.flags_i.N_1241\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__14582\,
            I => \N__14579\
        );

    \I__1792\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14574\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__14578\,
            I => \N__14570\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__14577\,
            I => \N__14564\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__14574\,
            I => \N__14561\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__14573\,
            I => \N__14556\
        );

    \I__1787\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14548\
        );

    \I__1786\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14548\
        );

    \I__1785\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14541\
        );

    \I__1784\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14541\
        );

    \I__1783\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14541\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__14561\,
            I => \N__14538\
        );

    \I__1781\ : InMux
    port map (
            O => \N__14560\,
            I => \N__14533\
        );

    \I__1780\ : InMux
    port map (
            O => \N__14559\,
            I => \N__14533\
        );

    \I__1779\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14530\
        );

    \I__1778\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14527\
        );

    \I__1777\ : InMux
    port map (
            O => \N__14554\,
            I => \N__14524\
        );

    \I__1776\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14521\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__14548\,
            I => \N__14516\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__14541\,
            I => \N__14516\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__14538\,
            I => \processor_zipi8.stack_pointer_0\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__14533\,
            I => \processor_zipi8.stack_pointer_0\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__14530\,
            I => \processor_zipi8.stack_pointer_0\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__14527\,
            I => \processor_zipi8.stack_pointer_0\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__14524\,
            I => \processor_zipi8.stack_pointer_0\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__14521\,
            I => \processor_zipi8.stack_pointer_0\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__14516\,
            I => \processor_zipi8.stack_pointer_0\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__14501\,
            I => \N__14498\
        );

    \I__1765\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__14495\,
            I => \N__14492\
        );

    \I__1763\ : Span4Mux_v
    port map (
            O => \N__14492\,
            I => \N__14488\
        );

    \I__1762\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14481\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__14488\,
            I => \N__14478\
        );

    \I__1760\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14473\
        );

    \I__1759\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14473\
        );

    \I__1758\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14468\
        );

    \I__1757\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14468\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__14481\,
            I => \N__14465\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__14478\,
            I => \processor_zipi8.stack_pointer_2\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__14473\,
            I => \processor_zipi8.stack_pointer_2\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__14468\,
            I => \processor_zipi8.stack_pointer_2\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__14465\,
            I => \processor_zipi8.stack_pointer_2\
        );

    \I__1751\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14449\
        );

    \I__1750\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14449\
        );

    \I__1749\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14446\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__14449\,
            I => \processor_zipi8.flags_i.N_54\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__14446\,
            I => \processor_zipi8.flags_i.N_54\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__14441\,
            I => \processor_zipi8.flags_i.m91_amZ0_cascade_\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__14438\,
            I => \processor_zipi8.flags_i.m25_ns_1_cascade_\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__14435\,
            I => \processor_zipi8.flags_i.N_26_0_cascade_\
        );

    \I__1743\ : InMux
    port map (
            O => \N__14432\,
            I => \N__14429\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__14429\,
            I => \processor_zipi8.flags_i.N_27_0\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__14426\,
            I => \processor_zipi8.flags_i.m20_ns_1_cascade_\
        );

    \I__1740\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14420\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__14420\,
            I => \processor_zipi8.flags_i.N_21_0\
        );

    \I__1738\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__14414\,
            I => \processor_zipi8.program_counter_i.half_pc_0_10\
        );

    \I__1736\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14408\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__14408\,
            I => \processor_zipi8.program_counter_i.un431_half_pc\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__14405\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_11_cascade_\
        );

    \I__1733\ : InMux
    port map (
            O => \N__14402\,
            I => \N__14399\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__14399\,
            I => \N__14395\
        );

    \I__1731\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__14395\,
            I => \processor_zipi8.address_11\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__14392\,
            I => \processor_zipi8.address_11\
        );

    \I__1728\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14384\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__14384\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_9\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__14381\,
            I => \N__14377\
        );

    \I__1725\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14374\
        );

    \I__1724\ : InMux
    port map (
            O => \N__14377\,
            I => \N__14371\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__14374\,
            I => \processor_zipi8.pc_vector_9\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__14371\,
            I => \processor_zipi8.pc_vector_9\
        );

    \I__1721\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14362\
        );

    \I__1720\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14359\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__14362\,
            I => \processor_zipi8.program_counter_i.carry_pc_52_8\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__14359\,
            I => \processor_zipi8.program_counter_i.carry_pc_52_8\
        );

    \I__1717\ : InMux
    port map (
            O => \N__14354\,
            I => \N__14350\
        );

    \I__1716\ : InMux
    port map (
            O => \N__14353\,
            I => \N__14347\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__14350\,
            I => \processor_zipi8.program_counter_i.carry_pc_58_9\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__14347\,
            I => \processor_zipi8.program_counter_i.carry_pc_58_9\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__14342\,
            I => \N__14339\
        );

    \I__1712\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14336\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__14336\,
            I => \processor_zipi8.flags_i.m49_ns_1\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__14333\,
            I => \processor_zipi8.flags_i.N_50_cascade_\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__14330\,
            I => \processor_zipi8.flags_i.N_51_cascade_\
        );

    \I__1708\ : InMux
    port map (
            O => \N__14327\,
            I => \N__14318\
        );

    \I__1707\ : InMux
    port map (
            O => \N__14326\,
            I => \N__14318\
        );

    \I__1706\ : InMux
    port map (
            O => \N__14325\,
            I => \N__14318\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__14318\,
            I => \processor_zipi8.flags_i.N_123_mux\
        );

    \I__1704\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14312\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__14312\,
            I => \processor_zipi8.flags_i.N_45\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__14309\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_4_cascade_\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__14306\,
            I => \processor_zipi8.program_counter_i.carry_pc_28_4_cascade_\
        );

    \I__1700\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14300\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__14300\,
            I => \processor_zipi8.program_counter_i.carry_pc_34_5\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__14297\,
            I => \N__14294\
        );

    \I__1697\ : InMux
    port map (
            O => \N__14294\,
            I => \N__14288\
        );

    \I__1696\ : InMux
    port map (
            O => \N__14293\,
            I => \N__14288\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__14288\,
            I => \N__14285\
        );

    \I__1694\ : Span4Mux_s2_h
    port map (
            O => \N__14285\,
            I => \N__14282\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__14282\,
            I => \processor_zipi8.pc_vector_6\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__14279\,
            I => \processor_zipi8.program_counter_i.carry_pc_34_5_cascade_\
        );

    \I__1691\ : InMux
    port map (
            O => \N__14276\,
            I => \N__14270\
        );

    \I__1690\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14270\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__14270\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_6\
        );

    \I__1688\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14264\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__14264\,
            I => \processor_zipi8.program_counter_i.carry_pc_40_6\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__14261\,
            I => \N__14257\
        );

    \I__1685\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14254\
        );

    \I__1684\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14251\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14245\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__14248\,
            I => \processor_zipi8.pc_vector_7\
        );

    \I__1680\ : Odrv12
    port map (
            O => \N__14245\,
            I => \processor_zipi8.pc_vector_7\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__14240\,
            I => \processor_zipi8.program_counter_i.carry_pc_40_6_cascade_\
        );

    \I__1678\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14233\
        );

    \I__1677\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14230\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__14233\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_7\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__14230\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_7\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__1673\ : CascadeBuf
    port map (
            O => \N__14222\,
            I => \N__14218\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__14221\,
            I => \N__14215\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__14218\,
            I => \N__14212\
        );

    \I__1670\ : CascadeBuf
    port map (
            O => \N__14215\,
            I => \N__14209\
        );

    \I__1669\ : CascadeBuf
    port map (
            O => \N__14212\,
            I => \N__14206\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__14209\,
            I => \N__14203\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__14206\,
            I => \N__14200\
        );

    \I__1666\ : CascadeBuf
    port map (
            O => \N__14203\,
            I => \N__14197\
        );

    \I__1665\ : CascadeBuf
    port map (
            O => \N__14200\,
            I => \N__14194\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__14197\,
            I => \N__14191\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__14194\,
            I => \N__14188\
        );

    \I__1662\ : CascadeBuf
    port map (
            O => \N__14191\,
            I => \N__14185\
        );

    \I__1661\ : CascadeBuf
    port map (
            O => \N__14188\,
            I => \N__14182\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__14185\,
            I => \N__14179\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__14182\,
            I => \N__14176\
        );

    \I__1658\ : CascadeBuf
    port map (
            O => \N__14179\,
            I => \N__14173\
        );

    \I__1657\ : CascadeBuf
    port map (
            O => \N__14176\,
            I => \N__14170\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__14173\,
            I => \N__14167\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__14170\,
            I => \N__14164\
        );

    \I__1654\ : CascadeBuf
    port map (
            O => \N__14167\,
            I => \N__14161\
        );

    \I__1653\ : CascadeBuf
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__14161\,
            I => \N__14155\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__14158\,
            I => \N__14152\
        );

    \I__1650\ : CascadeBuf
    port map (
            O => \N__14155\,
            I => \N__14149\
        );

    \I__1649\ : CascadeBuf
    port map (
            O => \N__14152\,
            I => \N__14146\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__14149\,
            I => \N__14143\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__14146\,
            I => \N__14140\
        );

    \I__1646\ : CascadeBuf
    port map (
            O => \N__14143\,
            I => \N__14137\
        );

    \I__1645\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14134\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__14137\,
            I => \N__14131\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__14134\,
            I => \N__14128\
        );

    \I__1642\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14125\
        );

    \I__1641\ : Span4Mux_s1_v
    port map (
            O => \N__14128\,
            I => \N__14116\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__14125\,
            I => \N__14116\
        );

    \I__1639\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14113\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__14123\,
            I => \N__14110\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__14122\,
            I => \N__14107\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__14121\,
            I => \N__14104\
        );

    \I__1635\ : Span4Mux_h
    port map (
            O => \N__14116\,
            I => \N__14101\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__14113\,
            I => \N__14098\
        );

    \I__1633\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14095\
        );

    \I__1632\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14092\
        );

    \I__1631\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14089\
        );

    \I__1630\ : Span4Mux_h
    port map (
            O => \N__14101\,
            I => \N__14086\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__14098\,
            I => address_7
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__14095\,
            I => address_7
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__14092\,
            I => address_7
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__14089\,
            I => address_7
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__14086\,
            I => address_7
        );

    \I__1624\ : InMux
    port map (
            O => \N__14075\,
            I => \N__14069\
        );

    \I__1623\ : InMux
    port map (
            O => \N__14074\,
            I => \N__14069\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__14069\,
            I => \N__14066\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__14066\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_5\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__1619\ : InMux
    port map (
            O => \N__14060\,
            I => \N__14054\
        );

    \I__1618\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14054\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__14054\,
            I => \N__14051\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__14051\,
            I => \processor_zipi8.pc_vector_5\
        );

    \I__1615\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14045\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__14045\,
            I => \processor_zipi8.program_counter_i.carry_pc_28_4\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__14042\,
            I => \N__14039\
        );

    \I__1612\ : CascadeBuf
    port map (
            O => \N__14039\,
            I => \N__14035\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__14038\,
            I => \N__14032\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__14035\,
            I => \N__14029\
        );

    \I__1609\ : CascadeBuf
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__1608\ : CascadeBuf
    port map (
            O => \N__14029\,
            I => \N__14023\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__14026\,
            I => \N__14020\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__14023\,
            I => \N__14017\
        );

    \I__1605\ : CascadeBuf
    port map (
            O => \N__14020\,
            I => \N__14014\
        );

    \I__1604\ : CascadeBuf
    port map (
            O => \N__14017\,
            I => \N__14011\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__14011\,
            I => \N__14005\
        );

    \I__1601\ : CascadeBuf
    port map (
            O => \N__14008\,
            I => \N__14002\
        );

    \I__1600\ : CascadeBuf
    port map (
            O => \N__14005\,
            I => \N__13999\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__14002\,
            I => \N__13996\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__13999\,
            I => \N__13993\
        );

    \I__1597\ : CascadeBuf
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__1596\ : CascadeBuf
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__13990\,
            I => \N__13984\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__13987\,
            I => \N__13981\
        );

    \I__1593\ : CascadeBuf
    port map (
            O => \N__13984\,
            I => \N__13978\
        );

    \I__1592\ : CascadeBuf
    port map (
            O => \N__13981\,
            I => \N__13975\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__13978\,
            I => \N__13972\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__1589\ : CascadeBuf
    port map (
            O => \N__13972\,
            I => \N__13966\
        );

    \I__1588\ : CascadeBuf
    port map (
            O => \N__13969\,
            I => \N__13963\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__13966\,
            I => \N__13960\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__13963\,
            I => \N__13957\
        );

    \I__1585\ : CascadeBuf
    port map (
            O => \N__13960\,
            I => \N__13954\
        );

    \I__1584\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__13954\,
            I => \N__13948\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__13951\,
            I => \N__13945\
        );

    \I__1581\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13942\
        );

    \I__1580\ : Span4Mux_s1_v
    port map (
            O => \N__13945\,
            I => \N__13933\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__13942\,
            I => \N__13933\
        );

    \I__1578\ : InMux
    port map (
            O => \N__13941\,
            I => \N__13930\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__13940\,
            I => \N__13927\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__13939\,
            I => \N__13924\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__13938\,
            I => \N__13921\
        );

    \I__1574\ : Span4Mux_h
    port map (
            O => \N__13933\,
            I => \N__13918\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__13930\,
            I => \N__13915\
        );

    \I__1572\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13912\
        );

    \I__1571\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13909\
        );

    \I__1570\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13906\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__13918\,
            I => \N__13903\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__13915\,
            I => address_5
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__13912\,
            I => address_5
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__13909\,
            I => address_5
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__13906\,
            I => address_5
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__13903\,
            I => address_5
        );

    \I__1563\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__13886\,
            I => \processor_zipi8.return_vector_11\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__13883\,
            I => \processor_zipi8.program_counter_i.un3_half_pcZ0_cascade_\
        );

    \I__1559\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13874\
        );

    \I__1558\ : InMux
    port map (
            O => \N__13879\,
            I => \N__13874\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__13874\,
            I => \processor_zipi8.flags_i.N_37\
        );

    \I__1556\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__13868\,
            I => \processor_zipi8.stack_memory_7\
        );

    \I__1554\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__13862\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_7\
        );

    \I__1552\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__13853\,
            I => \N__13850\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__13850\,
            I => \processor_zipi8.stack_memory_1\
        );

    \I__1548\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__13844\,
            I => \N__13841\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__13838\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_155\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__13835\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_195_cascade_\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__13832\,
            I => \N__13828\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__13831\,
            I => \N__13825\
        );

    \I__1541\ : CascadeBuf
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__1540\ : CascadeBuf
    port map (
            O => \N__13825\,
            I => \N__13819\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__13822\,
            I => \N__13816\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__13819\,
            I => \N__13813\
        );

    \I__1537\ : CascadeBuf
    port map (
            O => \N__13816\,
            I => \N__13810\
        );

    \I__1536\ : CascadeBuf
    port map (
            O => \N__13813\,
            I => \N__13807\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__13810\,
            I => \N__13804\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__13807\,
            I => \N__13801\
        );

    \I__1533\ : CascadeBuf
    port map (
            O => \N__13804\,
            I => \N__13798\
        );

    \I__1532\ : CascadeBuf
    port map (
            O => \N__13801\,
            I => \N__13795\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__13798\,
            I => \N__13792\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__13795\,
            I => \N__13789\
        );

    \I__1529\ : CascadeBuf
    port map (
            O => \N__13792\,
            I => \N__13786\
        );

    \I__1528\ : CascadeBuf
    port map (
            O => \N__13789\,
            I => \N__13783\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__13786\,
            I => \N__13780\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__13783\,
            I => \N__13777\
        );

    \I__1525\ : CascadeBuf
    port map (
            O => \N__13780\,
            I => \N__13774\
        );

    \I__1524\ : CascadeBuf
    port map (
            O => \N__13777\,
            I => \N__13771\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__13774\,
            I => \N__13768\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__13771\,
            I => \N__13765\
        );

    \I__1521\ : CascadeBuf
    port map (
            O => \N__13768\,
            I => \N__13762\
        );

    \I__1520\ : CascadeBuf
    port map (
            O => \N__13765\,
            I => \N__13759\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__13762\,
            I => \N__13756\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__13759\,
            I => \N__13753\
        );

    \I__1517\ : CascadeBuf
    port map (
            O => \N__13756\,
            I => \N__13750\
        );

    \I__1516\ : CascadeBuf
    port map (
            O => \N__13753\,
            I => \N__13747\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__13750\,
            I => \N__13744\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__13747\,
            I => \N__13741\
        );

    \I__1513\ : InMux
    port map (
            O => \N__13744\,
            I => \N__13737\
        );

    \I__1512\ : InMux
    port map (
            O => \N__13741\,
            I => \N__13734\
        );

    \I__1511\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13731\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__13737\,
            I => \N__13723\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__13734\,
            I => \N__13723\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__13731\,
            I => \N__13720\
        );

    \I__1507\ : InMux
    port map (
            O => \N__13730\,
            I => \N__13717\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__13729\,
            I => \N__13714\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__13728\,
            I => \N__13711\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__13723\,
            I => \N__13708\
        );

    \I__1503\ : Span4Mux_h
    port map (
            O => \N__13720\,
            I => \N__13705\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__13717\,
            I => \N__13702\
        );

    \I__1501\ : InMux
    port map (
            O => \N__13714\,
            I => \N__13699\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13711\,
            I => \N__13696\
        );

    \I__1499\ : Sp12to4
    port map (
            O => \N__13708\,
            I => \N__13693\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__13705\,
            I => address_6
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__13702\,
            I => address_6
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__13699\,
            I => address_6
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__13696\,
            I => address_6
        );

    \I__1494\ : Odrv12
    port map (
            O => \N__13693\,
            I => address_6
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__13682\,
            I => \N__13678\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__13681\,
            I => \N__13675\
        );

    \I__1491\ : CascadeBuf
    port map (
            O => \N__13678\,
            I => \N__13672\
        );

    \I__1490\ : CascadeBuf
    port map (
            O => \N__13675\,
            I => \N__13669\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__13672\,
            I => \N__13666\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__13669\,
            I => \N__13663\
        );

    \I__1487\ : CascadeBuf
    port map (
            O => \N__13666\,
            I => \N__13660\
        );

    \I__1486\ : CascadeBuf
    port map (
            O => \N__13663\,
            I => \N__13657\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__13660\,
            I => \N__13654\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__13657\,
            I => \N__13651\
        );

    \I__1483\ : CascadeBuf
    port map (
            O => \N__13654\,
            I => \N__13648\
        );

    \I__1482\ : CascadeBuf
    port map (
            O => \N__13651\,
            I => \N__13645\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__13648\,
            I => \N__13642\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__13645\,
            I => \N__13639\
        );

    \I__1479\ : CascadeBuf
    port map (
            O => \N__13642\,
            I => \N__13636\
        );

    \I__1478\ : CascadeBuf
    port map (
            O => \N__13639\,
            I => \N__13633\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__13636\,
            I => \N__13630\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__13633\,
            I => \N__13627\
        );

    \I__1475\ : CascadeBuf
    port map (
            O => \N__13630\,
            I => \N__13624\
        );

    \I__1474\ : CascadeBuf
    port map (
            O => \N__13627\,
            I => \N__13621\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__13624\,
            I => \N__13618\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__13621\,
            I => \N__13615\
        );

    \I__1471\ : CascadeBuf
    port map (
            O => \N__13618\,
            I => \N__13612\
        );

    \I__1470\ : CascadeBuf
    port map (
            O => \N__13615\,
            I => \N__13609\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__13612\,
            I => \N__13606\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__13609\,
            I => \N__13603\
        );

    \I__1467\ : CascadeBuf
    port map (
            O => \N__13606\,
            I => \N__13600\
        );

    \I__1466\ : CascadeBuf
    port map (
            O => \N__13603\,
            I => \N__13597\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__13600\,
            I => \N__13593\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__13597\,
            I => \N__13590\
        );

    \I__1463\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13587\
        );

    \I__1462\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13581\
        );

    \I__1461\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13578\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__13587\,
            I => \N__13575\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__13586\,
            I => \N__13572\
        );

    \I__1458\ : CascadeMux
    port map (
            O => \N__13585\,
            I => \N__13569\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__13584\,
            I => \N__13566\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__13581\,
            I => \N__13561\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__13578\,
            I => \N__13561\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__13575\,
            I => \N__13558\
        );

    \I__1453\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13555\
        );

    \I__1452\ : InMux
    port map (
            O => \N__13569\,
            I => \N__13552\
        );

    \I__1451\ : InMux
    port map (
            O => \N__13566\,
            I => \N__13549\
        );

    \I__1450\ : Span12Mux_s4_v
    port map (
            O => \N__13561\,
            I => \N__13546\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__13558\,
            I => address_4
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__13555\,
            I => address_4
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__13552\,
            I => address_4
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__13549\,
            I => address_4
        );

    \I__1445\ : Odrv12
    port map (
            O => \N__13546\,
            I => address_4
        );

    \I__1444\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13532\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__13532\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_4\
        );

    \I__1442\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13526\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__13526\,
            I => \N__13523\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__13523\,
            I => \processor_zipi8.stack_memory_6\
        );

    \I__1439\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13517\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__13517\,
            I => \N__13514\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__13514\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_6\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__13511\,
            I => \processor_zipi8.flags_i.N_125_mux_cascade_\
        );

    \I__1435\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__13505\,
            I => \processor_zipi8.stack_i.stack_bit\
        );

    \I__1433\ : InMux
    port map (
            O => \N__13502\,
            I => \N__13497\
        );

    \I__1432\ : InMux
    port map (
            O => \N__13501\,
            I => \N__13492\
        );

    \I__1431\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13492\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__13497\,
            I => \processor_zipi8.run\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__13492\,
            I => \processor_zipi8.run\
        );

    \I__1428\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13481\
        );

    \I__1427\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13481\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__13481\,
            I => \N__13478\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__1424\ : Span4Mux_h
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__1423\ : Span4Mux_h
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__13469\,
            I => \BTN1_c\
        );

    \I__1421\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__13463\,
            I => \processor_zipi8.stack_memory_2\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__13460\,
            I => \N__13456\
        );

    \I__1418\ : InMux
    port map (
            O => \N__13459\,
            I => \N__13451\
        );

    \I__1417\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13451\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__13451\,
            I => \processor_zipi8.special_bit\
        );

    \I__1415\ : IoInMux
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__1413\ : Span4Mux_s1_h
    port map (
            O => \N__13442\,
            I => \N__13439\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__13439\,
            I => \processor_zipi8.state_machine_i.bram_enable\
        );

    \I__1411\ : InMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__13433\,
            I => \processor_zipi8.stack_memory_11\
        );

    \I__1409\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13424\
        );

    \I__1408\ : InMux
    port map (
            O => \N__13429\,
            I => \N__13424\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__13424\,
            I => \N__13421\
        );

    \I__1406\ : Span4Mux_v
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__13418\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_6\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__13415\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_6_cascade_\
        );

    \I__1403\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13409\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__13409\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_6\
        );

    \I__1401\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13402\
        );

    \I__1400\ : InMux
    port map (
            O => \N__13405\,
            I => \N__13399\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__13402\,
            I => \N__13396\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__13399\,
            I => \N__13393\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__13396\,
            I => \N__13390\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__13393\,
            I => \N__13387\
        );

    \I__1395\ : Span4Mux_v
    port map (
            O => \N__13390\,
            I => \N__13384\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__13387\,
            I => \processor_zipi8.sy_6\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__13384\,
            I => \processor_zipi8.sy_6\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__13379\,
            I => \processor_zipi8.port_id_6_cascade_\
        );

    \I__1391\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__13373\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_6\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__13370\,
            I => \N__13367\
        );

    \I__1388\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13363\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__13366\,
            I => \N__13359\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__13363\,
            I => \N__13356\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__13362\,
            I => \N__13352\
        );

    \I__1384\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13348\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__13356\,
            I => \N__13345\
        );

    \I__1382\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13338\
        );

    \I__1381\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13338\
        );

    \I__1380\ : InMux
    port map (
            O => \N__13351\,
            I => \N__13338\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__13348\,
            I => \processor_zipi8.port_id_6\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__13345\,
            I => \processor_zipi8.port_id_6\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__13338\,
            I => \processor_zipi8.port_id_6\
        );

    \I__1376\ : InMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__13328\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_6\
        );

    \I__1374\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13319\
        );

    \I__1373\ : InMux
    port map (
            O => \N__13324\,
            I => \N__13319\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__13319\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_5\
        );

    \I__1371\ : InMux
    port map (
            O => \N__13316\,
            I => \N__13312\
        );

    \I__1370\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13309\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__13312\,
            I => \N__13304\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13304\
        );

    \I__1367\ : Odrv12
    port map (
            O => \N__13304\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_6\
        );

    \I__1366\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13295\
        );

    \I__1365\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13295\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__13295\,
            I => \N__13292\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__13292\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_7\
        );

    \I__1362\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__13286\,
            I => \processor_zipi8.spm_data_5\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__13283\,
            I => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202_cascade_\
        );

    \I__1359\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13274\
        );

    \I__1358\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13274\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__13274\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_5\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__1355\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13265\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__13265\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_5\
        );

    \I__1353\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13256\
        );

    \I__1352\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13256\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13253\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__13253\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_6\
        );

    \I__1349\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13247\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__1347\ : Span4Mux_s2_h
    port map (
            O => \N__13244\,
            I => \N__13240\
        );

    \I__1346\ : InMux
    port map (
            O => \N__13243\,
            I => \N__13237\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__13240\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__13237\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7\
        );

    \I__1343\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__13226\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_7\
        );

    \I__1340\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13217\
        );

    \I__1339\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13217\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__13214\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_5\
        );

    \I__1336\ : InMux
    port map (
            O => \N__13211\,
            I => \N__13205\
        );

    \I__1335\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13205\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__13205\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_6\
        );

    \I__1333\ : InMux
    port map (
            O => \N__13202\,
            I => \N__13198\
        );

    \I__1332\ : InMux
    port map (
            O => \N__13201\,
            I => \N__13195\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__13198\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__13195\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__13190\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_6_cascade_\
        );

    \I__1328\ : InMux
    port map (
            O => \N__13187\,
            I => \N__13184\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__13184\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_6\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__13181\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_6_cascade_\
        );

    \I__1325\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13172\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__13172\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_6\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__13169\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_6_cascade_\
        );

    \I__1321\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13163\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__13163\,
            I => \N__13160\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__13160\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_6\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__13157\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_6_cascade_\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__13154\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_6_cascade_\
        );

    \I__1316\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13147\
        );

    \I__1315\ : InMux
    port map (
            O => \N__13150\,
            I => \N__13144\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__13147\,
            I => \N__13139\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__13144\,
            I => \N__13139\
        );

    \I__1312\ : Span4Mux_v
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__13136\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_7\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__13133\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_6_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__13130\,
            I => \N__13126\
        );

    \I__1308\ : InMux
    port map (
            O => \N__13129\,
            I => \N__13123\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__13126\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__13123\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__13118\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_7_cascade_\
        );

    \I__1304\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13112\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__13112\,
            I => \N__13109\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__13109\,
            I => \N__13106\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__13106\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIK2TR1_7\
        );

    \I__1300\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13099\
        );

    \I__1299\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13096\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__13099\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__13096\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7\
        );

    \I__1296\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13088\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__13088\,
            I => \processor_zipi8.alu_result_3\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__13085\,
            I => \processor_zipi8.flags_i.m82_1_cascade_\
        );

    \I__1293\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13079\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__13079\,
            I => \processor_zipi8.flags_i.m82_1\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__13076\,
            I => \N__13073\
        );

    \I__1290\ : InMux
    port map (
            O => \N__13073\,
            I => \N__13070\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__13070\,
            I => \N__13067\
        );

    \I__1288\ : Span4Mux_h
    port map (
            O => \N__13067\,
            I => \N__13064\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__13064\,
            I => \N__13061\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__13061\,
            I => \processor_zipi8.zero_flag_RNIJSPM4\
        );

    \I__1285\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13055\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__13055\,
            I => \processor_zipi8.flags_i.N_55\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__13052\,
            I => \processor_zipi8.flags_i.m61_ns_1_cascade_\
        );

    \I__1282\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13046\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__13046\,
            I => \N__13043\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__13043\,
            I => \processor_zipi8.pc_vector_8\
        );

    \I__1279\ : CascadeMux
    port map (
            O => \N__13040\,
            I => \processor_zipi8.program_counter_i.carry_pc_46_7_cascade_\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__13037\,
            I => \N__13033\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__13036\,
            I => \N__13030\
        );

    \I__1276\ : CascadeBuf
    port map (
            O => \N__13033\,
            I => \N__13027\
        );

    \I__1275\ : CascadeBuf
    port map (
            O => \N__13030\,
            I => \N__13024\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__13027\,
            I => \N__13021\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__13024\,
            I => \N__13018\
        );

    \I__1272\ : CascadeBuf
    port map (
            O => \N__13021\,
            I => \N__13015\
        );

    \I__1271\ : CascadeBuf
    port map (
            O => \N__13018\,
            I => \N__13012\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__13015\,
            I => \N__13009\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__13012\,
            I => \N__13006\
        );

    \I__1268\ : CascadeBuf
    port map (
            O => \N__13009\,
            I => \N__13003\
        );

    \I__1267\ : CascadeBuf
    port map (
            O => \N__13006\,
            I => \N__13000\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__13003\,
            I => \N__12997\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__13000\,
            I => \N__12994\
        );

    \I__1264\ : CascadeBuf
    port map (
            O => \N__12997\,
            I => \N__12991\
        );

    \I__1263\ : CascadeBuf
    port map (
            O => \N__12994\,
            I => \N__12988\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__12991\,
            I => \N__12985\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__12988\,
            I => \N__12982\
        );

    \I__1260\ : CascadeBuf
    port map (
            O => \N__12985\,
            I => \N__12979\
        );

    \I__1259\ : CascadeBuf
    port map (
            O => \N__12982\,
            I => \N__12976\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__12979\,
            I => \N__12973\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__12976\,
            I => \N__12970\
        );

    \I__1256\ : CascadeBuf
    port map (
            O => \N__12973\,
            I => \N__12967\
        );

    \I__1255\ : CascadeBuf
    port map (
            O => \N__12970\,
            I => \N__12964\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__12967\,
            I => \N__12961\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__12964\,
            I => \N__12958\
        );

    \I__1252\ : CascadeBuf
    port map (
            O => \N__12961\,
            I => \N__12955\
        );

    \I__1251\ : CascadeBuf
    port map (
            O => \N__12958\,
            I => \N__12952\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__12955\,
            I => \N__12948\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__12952\,
            I => \N__12945\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__12951\,
            I => \N__12940\
        );

    \I__1247\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12936\
        );

    \I__1246\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12933\
        );

    \I__1245\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12930\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__12943\,
            I => \N__12927\
        );

    \I__1243\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12924\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__12939\,
            I => \N__12921\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__12936\,
            I => \N__12918\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__12933\,
            I => \N__12915\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__12930\,
            I => \N__12912\
        );

    \I__1238\ : InMux
    port map (
            O => \N__12927\,
            I => \N__12909\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__12924\,
            I => \N__12906\
        );

    \I__1236\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12903\
        );

    \I__1235\ : Span4Mux_v
    port map (
            O => \N__12918\,
            I => \N__12898\
        );

    \I__1234\ : Span4Mux_v
    port map (
            O => \N__12915\,
            I => \N__12898\
        );

    \I__1233\ : Span4Mux_h
    port map (
            O => \N__12912\,
            I => \N__12895\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__12909\,
            I => \N__12890\
        );

    \I__1231\ : Span4Mux_h
    port map (
            O => \N__12906\,
            I => \N__12890\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__12903\,
            I => \N__12885\
        );

    \I__1229\ : Sp12to4
    port map (
            O => \N__12898\,
            I => \N__12885\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__12895\,
            I => address_8
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__12890\,
            I => address_8
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__12885\,
            I => address_8
        );

    \I__1225\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__12875\,
            I => \N__12871\
        );

    \I__1223\ : InMux
    port map (
            O => \N__12874\,
            I => \N__12868\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__12871\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_8\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__12868\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_8\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__12863\,
            I => \processor_zipi8.flags_i.zero_flag_3_cascade_\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__12860\,
            I => \N__12857\
        );

    \I__1218\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__12854\,
            I => \processor_zipi8.shadow_zero_flag\
        );

    \I__1216\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__12848\,
            I => \N__12845\
        );

    \I__1214\ : Span12Mux_s3_v
    port map (
            O => \N__12845\,
            I => \N__12842\
        );

    \I__1213\ : Odrv12
    port map (
            O => \N__12842\,
            I => \processor_zipi8.alu_result_7\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__12839\,
            I => \processor_zipi8.alu_result_6_cascade_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__12833\,
            I => \processor_zipi8.flags_i.zero_flag_3_0_5\
        );

    \I__1209\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12827\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__12827\,
            I => \processor_zipi8.alu_result_5\
        );

    \I__1207\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12821\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__12821\,
            I => \N__12818\
        );

    \I__1205\ : Span4Mux_s3_v
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__1204\ : Span4Mux_v
    port map (
            O => \N__12815\,
            I => \N__12812\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__12812\,
            I => \processor_zipi8.stack_i.stack_zero_flag\
        );

    \I__1202\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__12806\,
            I => \processor_zipi8.stack_i.shadow_zero_value\
        );

    \I__1200\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__12800\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_8\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__12797\,
            I => \processor_zipi8.pc_vector_8_cascade_\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__12794\,
            I => \processor_zipi8.program_counter_i.half_pc_0_0_9_cascade_\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__12791\,
            I => \N__12787\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__12790\,
            I => \N__12784\
        );

    \I__1194\ : CascadeBuf
    port map (
            O => \N__12787\,
            I => \N__12781\
        );

    \I__1193\ : CascadeBuf
    port map (
            O => \N__12784\,
            I => \N__12778\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__12781\,
            I => \N__12775\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__12778\,
            I => \N__12772\
        );

    \I__1190\ : CascadeBuf
    port map (
            O => \N__12775\,
            I => \N__12769\
        );

    \I__1189\ : CascadeBuf
    port map (
            O => \N__12772\,
            I => \N__12766\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__12769\,
            I => \N__12763\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__12766\,
            I => \N__12760\
        );

    \I__1186\ : CascadeBuf
    port map (
            O => \N__12763\,
            I => \N__12757\
        );

    \I__1185\ : CascadeBuf
    port map (
            O => \N__12760\,
            I => \N__12754\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__12757\,
            I => \N__12751\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__12754\,
            I => \N__12748\
        );

    \I__1182\ : CascadeBuf
    port map (
            O => \N__12751\,
            I => \N__12745\
        );

    \I__1181\ : CascadeBuf
    port map (
            O => \N__12748\,
            I => \N__12742\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__12745\,
            I => \N__12739\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__12742\,
            I => \N__12736\
        );

    \I__1178\ : CascadeBuf
    port map (
            O => \N__12739\,
            I => \N__12733\
        );

    \I__1177\ : CascadeBuf
    port map (
            O => \N__12736\,
            I => \N__12730\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__12733\,
            I => \N__12727\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__12730\,
            I => \N__12724\
        );

    \I__1174\ : CascadeBuf
    port map (
            O => \N__12727\,
            I => \N__12721\
        );

    \I__1173\ : CascadeBuf
    port map (
            O => \N__12724\,
            I => \N__12718\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__12721\,
            I => \N__12715\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__12718\,
            I => \N__12712\
        );

    \I__1170\ : CascadeBuf
    port map (
            O => \N__12715\,
            I => \N__12709\
        );

    \I__1169\ : CascadeBuf
    port map (
            O => \N__12712\,
            I => \N__12706\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__12709\,
            I => \N__12703\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__12706\,
            I => \N__12700\
        );

    \I__1166\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12696\
        );

    \I__1165\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12693\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__12699\,
            I => \N__12688\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__12696\,
            I => \N__12685\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__12693\,
            I => \N__12682\
        );

    \I__1161\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12679\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__12691\,
            I => \N__12675\
        );

    \I__1159\ : InMux
    port map (
            O => \N__12688\,
            I => \N__12672\
        );

    \I__1158\ : Span4Mux_s1_v
    port map (
            O => \N__12685\,
            I => \N__12667\
        );

    \I__1157\ : Span4Mux_s2_h
    port map (
            O => \N__12682\,
            I => \N__12667\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__12679\,
            I => \N__12664\
        );

    \I__1155\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12661\
        );

    \I__1154\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12658\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__12672\,
            I => \N__12655\
        );

    \I__1152\ : Span4Mux_h
    port map (
            O => \N__12667\,
            I => \N__12652\
        );

    \I__1151\ : Span4Mux_v
    port map (
            O => \N__12664\,
            I => \N__12645\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__12661\,
            I => \N__12645\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__12658\,
            I => \N__12645\
        );

    \I__1148\ : Span4Mux_h
    port map (
            O => \N__12655\,
            I => \N__12640\
        );

    \I__1147\ : Span4Mux_h
    port map (
            O => \N__12652\,
            I => \N__12640\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__12645\,
            I => address_9
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__12640\,
            I => address_9
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__12635\,
            I => \processor_zipi8.program_counter_i.un380_half_pc_cascade_\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__12632\,
            I => \processor_zipi8.program_counter_i.half_pc_0_10_cascade_\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__12629\,
            I => \N__12625\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__12628\,
            I => \N__12622\
        );

    \I__1140\ : CascadeBuf
    port map (
            O => \N__12625\,
            I => \N__12619\
        );

    \I__1139\ : CascadeBuf
    port map (
            O => \N__12622\,
            I => \N__12616\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__12619\,
            I => \N__12613\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__12616\,
            I => \N__12610\
        );

    \I__1136\ : CascadeBuf
    port map (
            O => \N__12613\,
            I => \N__12607\
        );

    \I__1135\ : CascadeBuf
    port map (
            O => \N__12610\,
            I => \N__12604\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__12607\,
            I => \N__12601\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__12604\,
            I => \N__12598\
        );

    \I__1132\ : CascadeBuf
    port map (
            O => \N__12601\,
            I => \N__12595\
        );

    \I__1131\ : CascadeBuf
    port map (
            O => \N__12598\,
            I => \N__12592\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__12595\,
            I => \N__12589\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__12592\,
            I => \N__12586\
        );

    \I__1128\ : CascadeBuf
    port map (
            O => \N__12589\,
            I => \N__12583\
        );

    \I__1127\ : CascadeBuf
    port map (
            O => \N__12586\,
            I => \N__12580\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__12583\,
            I => \N__12577\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__12580\,
            I => \N__12574\
        );

    \I__1124\ : CascadeBuf
    port map (
            O => \N__12577\,
            I => \N__12571\
        );

    \I__1123\ : CascadeBuf
    port map (
            O => \N__12574\,
            I => \N__12568\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__12571\,
            I => \N__12565\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__12568\,
            I => \N__12562\
        );

    \I__1120\ : CascadeBuf
    port map (
            O => \N__12565\,
            I => \N__12559\
        );

    \I__1119\ : CascadeBuf
    port map (
            O => \N__12562\,
            I => \N__12556\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__12559\,
            I => \N__12553\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__12556\,
            I => \N__12550\
        );

    \I__1116\ : CascadeBuf
    port map (
            O => \N__12553\,
            I => \N__12547\
        );

    \I__1115\ : CascadeBuf
    port map (
            O => \N__12550\,
            I => \N__12544\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__12547\,
            I => \N__12540\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__12544\,
            I => \N__12537\
        );

    \I__1112\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12533\
        );

    \I__1111\ : InMux
    port map (
            O => \N__12540\,
            I => \N__12529\
        );

    \I__1110\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12526\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__12536\,
            I => \N__12523\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__12533\,
            I => \N__12520\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__12532\,
            I => \N__12517\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__12529\,
            I => \N__12512\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__12526\,
            I => \N__12512\
        );

    \I__1104\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12509\
        );

    \I__1103\ : Span4Mux_v
    port map (
            O => \N__12520\,
            I => \N__12506\
        );

    \I__1102\ : InMux
    port map (
            O => \N__12517\,
            I => \N__12503\
        );

    \I__1101\ : Span4Mux_s3_v
    port map (
            O => \N__12512\,
            I => \N__12500\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__12509\,
            I => \N__12495\
        );

    \I__1099\ : Sp12to4
    port map (
            O => \N__12506\,
            I => \N__12490\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__12503\,
            I => \N__12490\
        );

    \I__1097\ : Span4Mux_h
    port map (
            O => \N__12500\,
            I => \N__12487\
        );

    \I__1096\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12482\
        );

    \I__1095\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12482\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__12495\,
            I => \N__12479\
        );

    \I__1093\ : Span12Mux_s11_h
    port map (
            O => \N__12490\,
            I => \N__12476\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__12487\,
            I => \N__12473\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__12482\,
            I => address_10
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__12479\,
            I => address_10
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__12476\,
            I => address_10
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__12473\,
            I => address_10
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__12464\,
            I => \N__12461\
        );

    \I__1086\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__12458\,
            I => \N__12455\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__12455\,
            I => \N__12452\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__12452\,
            I => \processor_zipi8.return_vector_10\
        );

    \I__1082\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12446\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__12446\,
            I => \processor_zipi8.program_counter_i.un395_half_pcZ0\
        );

    \I__1080\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12440\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__12440\,
            I => \processor_zipi8.program_counter_i.carry_pc_46_7\
        );

    \I__1078\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12434\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__12431\,
            I => \processor_zipi8.stack_memory_9\
        );

    \I__1075\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12425\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__12425\,
            I => \N__12422\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__12422\,
            I => \processor_zipi8.stack_memory_4\
        );

    \I__1072\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__12413\,
            I => \N__12410\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__12410\,
            I => \processor_zipi8.stack_memory_8\
        );

    \I__1068\ : InMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__12404\,
            I => \N__12401\
        );

    \I__1066\ : Span4Mux_v
    port map (
            O => \N__12401\,
            I => \N__12398\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__12398\,
            I => \processor_zipi8.stack_memory_10\
        );

    \I__1064\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__1062\ : Span4Mux_h
    port map (
            O => \N__12389\,
            I => \N__12386\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__12386\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_9\
        );

    \I__1060\ : InMux
    port map (
            O => \N__12383\,
            I => \N__12379\
        );

    \I__1059\ : InMux
    port map (
            O => \N__12382\,
            I => \N__12376\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__12379\,
            I => \N__12371\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__12376\,
            I => \N__12371\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__12371\,
            I => \processor_zipi8.sy_5\
        );

    \I__1055\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12364\
        );

    \I__1054\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12361\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__12364\,
            I => \N__12358\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__12361\,
            I => \N__12355\
        );

    \I__1051\ : Span4Mux_h
    port map (
            O => \N__12358\,
            I => \N__12350\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__12355\,
            I => \N__12350\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__12350\,
            I => \processor_zipi8.sy_7\
        );

    \I__1048\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12344\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__12344\,
            I => \N__12341\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__12341\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_7\
        );

    \I__1045\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12335\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__12335\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_7\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__12332\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_7_cascade_\
        );

    \I__1042\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12326\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__12326\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_7\
        );

    \I__1040\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12320\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__12320\,
            I => \N__12317\
        );

    \I__1038\ : Span4Mux_v
    port map (
            O => \N__12317\,
            I => \N__12314\
        );

    \I__1037\ : Span4Mux_s1_h
    port map (
            O => \N__12314\,
            I => \N__12311\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__12311\,
            I => \processor_zipi8.stack_memory_5\
        );

    \I__1035\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12305\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__12305\,
            I => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_5\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__12302\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_5_cascade_\
        );

    \I__1032\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12296\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__12296\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_5\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__12293\,
            I => \processor_zipi8.port_id_5_cascade_\
        );

    \I__1029\ : InMux
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__12287\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_5\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__12284\,
            I => \N__12280\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__12283\,
            I => \N__12277\
        );

    \I__1025\ : InMux
    port map (
            O => \N__12280\,
            I => \N__12274\
        );

    \I__1024\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12271\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__12274\,
            I => \N__12268\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__12271\,
            I => \N__12265\
        );

    \I__1021\ : Span4Mux_v
    port map (
            O => \N__12268\,
            I => \N__12259\
        );

    \I__1020\ : Span4Mux_h
    port map (
            O => \N__12265\,
            I => \N__12256\
        );

    \I__1019\ : InMux
    port map (
            O => \N__12264\,
            I => \N__12249\
        );

    \I__1018\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12249\
        );

    \I__1017\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12249\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__12259\,
            I => \processor_zipi8.port_id_5\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__12256\,
            I => \processor_zipi8.port_id_5\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__12249\,
            I => \processor_zipi8.port_id_5\
        );

    \I__1013\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__12239\,
            I => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_5\
        );

    \I__1011\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12233\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__12230\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI88F42_7\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__12227\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV3DI8_7_cascade_\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__12224\,
            I => \N__12221\
        );

    \I__1006\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12218\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__1004\ : Odrv12
    port map (
            O => \N__12215\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIM5NP1_7\
        );

    \I__1003\ : InMux
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__12209\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_7\
        );

    \I__1001\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__12203\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINR4G8_7\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__12200\,
            I => \processor_zipi8.port_id_7_cascade_\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__12197\,
            I => \N__12193\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__12196\,
            I => \N__12190\
        );

    \I__996\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12187\
        );

    \I__995\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12184\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12181\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__12181\,
            I => \N__12172\
        );

    \I__991\ : Span4Mux_h
    port map (
            O => \N__12178\,
            I => \N__12169\
        );

    \I__990\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12162\
        );

    \I__989\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12162\
        );

    \I__988\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12162\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__12172\,
            I => \processor_zipi8.port_id_7\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__12169\,
            I => \processor_zipi8.port_id_7\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__12162\,
            I => \processor_zipi8.port_id_7\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__12155\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_5_cascade_\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__12152\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_5_cascade_\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__12149\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_5_cascade_\
        );

    \I__981\ : InMux
    port map (
            O => \N__12146\,
            I => \N__12143\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__12143\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_5\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__12140\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_5_cascade_\
        );

    \I__978\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__12134\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_5\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__12131\,
            I => \processor_zipi8.flags_i.un5_shift_carry_value_cascade_\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__12128\,
            I => \processor_zipi8.flags_i.shift_carry_value_1_0_0_cascade_\
        );

    \I__974\ : InMux
    port map (
            O => \N__12125\,
            I => \N__12122\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__12122\,
            I => \N__12119\
        );

    \I__972\ : Span4Mux_v
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__12116\,
            I => \processor_zipi8.stack_i.data_out_ram_0\
        );

    \I__970\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12110\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__12110\,
            I => \processor_zipi8.shadow_carry_flag\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__12107\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_7_cascade_\
        );

    \I__967\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12098\
        );

    \I__966\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12098\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__12098\,
            I => \N__12095\
        );

    \I__964\ : Span4Mux_v
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__12092\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_7\
        );

    \I__962\ : InMux
    port map (
            O => \N__12089\,
            I => \N__12086\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__12086\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_7\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__12083\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_7_cascade_\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__12080\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_7_cascade_\
        );

    \I__958\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__12074\,
            I => \N__12071\
        );

    \I__956\ : Span4Mux_s1_h
    port map (
            O => \N__12071\,
            I => \N__12068\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__12068\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_7\
        );

    \I__954\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__12062\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_7\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__12059\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_7_cascade_\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__12056\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_7_cascade_\
        );

    \I__950\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12050\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__12050\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_7\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__12047\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_7_cascade_\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__12044\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_7_cascade_\
        );

    \I__946\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12035\
        );

    \I__945\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12035\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__12035\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_7\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__12032\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_7_cascade_\
        );

    \I__942\ : InMux
    port map (
            O => \N__12029\,
            I => \N__12023\
        );

    \I__941\ : InMux
    port map (
            O => \N__12028\,
            I => \N__12023\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__12023\,
            I => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_7\
        );

    \processor_zipi8.state_machine_i.t_state_RNIA073_2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__13448\,
            GLOBALBUFFEROUTPUT => bram_enable_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__7_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__33312\,
            in1 => \N__32974\,
            in2 => \N__36522\,
            in3 => \N__34765\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33634\,
            ce => \N__14864\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_7_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37469\,
            in1 => \N__16426\,
            in2 => \_gnd_net_\,
            in3 => \N__13102\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__6_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34084\,
            in1 => \N__29265\,
            in2 => \N__36701\,
            in3 => \N__29707\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33623\,
            ce => \N__25944\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__7_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__32973\,
            in1 => \N__34085\,
            in2 => \N__36700\,
            in3 => \N__33340\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33623\,
            ce => \N__25944\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_7_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34079\,
            in1 => \N__32824\,
            in2 => \N__33320\,
            in3 => \N__36050\,
            lcout => \processor_zipi8.alu_result_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__7_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36051\,
            in1 => \N__33270\,
            in2 => \N__32898\,
            in3 => \N__34080\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33614\,
            ce => \N__25339\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_7_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12028\,
            in1 => \N__13150\,
            in2 => \_gnd_net_\,
            in3 => \N__37498\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_7_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37499\,
            in1 => \N__23782\,
            in2 => \_gnd_net_\,
            in3 => \N__12040\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_7_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__12053\,
            in1 => \N__28653\,
            in2 => \N__12047\,
            in3 => \N__29013\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_7_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28654\,
            in1 => \N__20411\,
            in2 => \N__12044\,
            in3 => \N__20453\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIP1UE1_7_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__12041\,
            in1 => \N__31699\,
            in2 => \N__23786\,
            in3 => \N__30993\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI88F42_7_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31700\,
            in1 => \N__13151\,
            in2 => \N__12032\,
            in3 => \N__12029\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI88F42_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_7_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13300\,
            in1 => \N__12103\,
            in2 => \_gnd_net_\,
            in3 => \N__37496\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI92021_7_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__13202\,
            in1 => \N__31702\,
            in2 => \N__31016\,
            in3 => \N__16469\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIM5NP1_7_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__13301\,
            in1 => \N__31750\,
            in2 => \N__12107\,
            in3 => \N__12104\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIM5NP1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_7_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37497\,
            in1 => \N__16468\,
            in2 => \_gnd_net_\,
            in3 => \N__13201\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_7_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__29005\,
            in1 => \N__12089\,
            in2 => \N__12083\,
            in3 => \N__28655\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_7_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28656\,
            in1 => \N__13232\,
            in2 => \N__12080\,
            in3 => \N__12077\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_7_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__12065\,
            in1 => \N__25669\,
            in2 => \N__12059\,
            in3 => \N__25792\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_7_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25670\,
            in1 => \N__28310\,
            in2 => \N__12056\,
            in3 => \N__20933\,
            lcout => \processor_zipi8.sy_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_5_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13324\,
            in1 => \N__13279\,
            in2 => \_gnd_net_\,
            in3 => \N__37494\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI5UV11_5_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__13223\,
            in1 => \N__31696\,
            in2 => \N__31015\,
            in3 => \N__16496\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIETMP1_5_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__13325\,
            in1 => \N__31697\,
            in2 => \N__12155\,
            in3 => \N__13280\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_5_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__18104\,
            in1 => \N__12137\,
            in2 => \N__13271\,
            in3 => \N__28622\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_5_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__24986\,
            in1 => \N__25660\,
            in2 => \N__12152\,
            in3 => \N__25761\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_5_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25661\,
            in1 => \N__22697\,
            in2 => \N__12149\,
            in3 => \N__20399\,
            lcout => \processor_zipi8.sy_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_5_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16495\,
            in1 => \N__13222\,
            in2 => \_gnd_net_\,
            in3 => \N__37495\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_5_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__12146\,
            in1 => \N__28621\,
            in2 => \N__12140\,
            in3 => \N__29004\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.shift_carry_RNO_1_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__16679\,
            in1 => \N__17102\,
            in2 => \_gnd_net_\,
            in3 => \N__24316\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.un5_shift_carry_value_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.shift_carry_RNO_0_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000111"
        )
    port map (
            in0 => \N__25783\,
            in1 => \N__24318\,
            in2 => \N__12131\,
            in3 => \N__12113\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.shift_carry_value_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.shift_carry_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__17121\,
            in1 => \N__24317\,
            in2 => \N__12128\,
            in3 => \N__21113\,
            lcout => \processor_zipi8.flags_i.shift_carryZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.shadow_carry_flag_0_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12125\,
            lcout => \processor_zipi8.shadow_carry_flag\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU7BG4_7_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__12236\,
            in1 => \N__27439\,
            in2 => \N__20252\,
            in3 => \N__27636\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV3DI8_7_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__27441\,
            in1 => \N__28259\,
            in2 => \N__22883\,
            in3 => \N__20222\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV3DI8_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5S0IH_7_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__12206\,
            in1 => \_gnd_net_\,
            in2 => \N__12227\,
            in3 => \N__22233\,
            lcout => \processor_zipi8.sx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINR4G8_7_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__27440\,
            in1 => \N__13115\,
            in2 => \N__12224\,
            in3 => \N__12212\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINR4G8_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_7_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111110111"
        )
    port map (
            in0 => \N__12176\,
            in1 => \N__19588\,
            in2 => \N__16684\,
            in3 => \N__19639\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12368\,
            in1 => \N__21447\,
            in2 => \_gnd_net_\,
            in3 => \N__25782\,
            lcout => \processor_zipi8.port_id_7\,
            ltout => \processor_zipi8.port_id_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_7_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__16667\,
            in1 => \N__19208\,
            in2 => \N__12200\,
            in3 => \N__19589\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_7_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110111"
        )
    port map (
            in0 => \N__19207\,
            in1 => \N__12177\,
            in2 => \N__16683\,
            in3 => \N__24013\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_7_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__12175\,
            in1 => \N__19486\,
            in2 => \N__16685\,
            in3 => \N__19799\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_7_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12347\,
            in1 => \N__12338\,
            in2 => \N__12332\,
            in3 => \N__12329\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_5_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNID2G21_5_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29015\,
            in1 => \N__12308\,
            in2 => \_gnd_net_\,
            in3 => \N__21446\,
            lcout => \processor_zipi8.pc_vector_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_5_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__12262\,
            in1 => \N__19478\,
            in2 => \N__18784\,
            in3 => \N__19797\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_5_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__12242\,
            in1 => \N__12290\,
            in2 => \N__12302\,
            in3 => \N__12299\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_5_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__12263\,
            in1 => \N__19580\,
            in2 => \N__18783\,
            in3 => \N__19201\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_2_0_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12383\,
            in1 => \N__21452\,
            in2 => \_gnd_net_\,
            in3 => \N__29014\,
            lcout => \processor_zipi8.port_id_5\,
            ltout => \processor_zipi8.port_id_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_5_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__18765\,
            in1 => \N__19579\,
            in2 => \N__12293\,
            in3 => \N__19632\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_5_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000111"
        )
    port map (
            in0 => \N__19200\,
            in1 => \N__12264\,
            in2 => \N__24014\,
            in3 => \N__18766\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_9_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12437\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_4_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12428\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIG4G21_7_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13865\,
            in1 => \N__21453\,
            in2 => \_gnd_net_\,
            in3 => \N__25784\,
            lcout => \processor_zipi8.pc_vector_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_8_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12419\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_10_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12407\,
            lcout => \processor_zipi8.return_vector_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIJ6G21_9_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12395\,
            in1 => \N__21455\,
            in2 => \_gnd_net_\,
            in3 => \N__31694\,
            lcout => \processor_zipi8.pc_vector_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNING29O_5_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__12382\,
            in1 => \N__17882\,
            in2 => \N__13940\,
            in3 => \N__17800\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIOI39O_6_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__17801\,
            in1 => \N__13730\,
            in2 => \N__17890\,
            in3 => \N__13406\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIPK49O_7_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__12367\,
            in1 => \N__17886\,
            in2 => \N__14123\,
            in3 => \N__17802\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNII5G21_8_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12803\,
            in1 => \N__21454\,
            in2 => \_gnd_net_\,
            in3 => \N__31021\,
            lcout => \processor_zipi8.pc_vector_8\,
            ltout => \processor_zipi8.pc_vector_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_8_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100110011001"
        )
    port map (
            in0 => \N__12878\,
            in1 => \N__12443\,
            in2 => \N__12797\,
            in3 => \N__15939\,
            lcout => address_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33622\,
            ce => \N__15763\,
            sr => \N__17401\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNI9LLGO_9_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__17803\,
            in1 => \N__12678\,
            in2 => \N__17891\,
            in3 => \N__21706\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_9\,
            ltout => \processor_zipi8.program_counter_i.half_pc_0_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_9_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000010001111"
        )
    port map (
            in0 => \N__14380\,
            in1 => \N__15940\,
            in2 => \N__12794\,
            in3 => \N__14366\,
            lcout => address_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33622\,
            ce => \N__15763\,
            sr => \N__17401\
        );

    \processor_zipi8.program_counter_i.pc_RNIDL1F5_10_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12498\,
            lcout => OPEN,
            ltout => \processor_zipi8.program_counter_i.un380_half_pc_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_RNIDJA501_10_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__17861\,
            in1 => \N__22013\,
            in2 => \N__12635\,
            in3 => \N__12449\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_10\,
            ltout => \processor_zipi8.program_counter_i.half_pc_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_10_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__19058\,
            in1 => \N__12499\,
            in2 => \N__12632\,
            in3 => \N__14354\,
            lcout => address_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33626\,
            ce => 'H',
            sr => \N__17429\
        );

    \processor_zipi8.program_counter_i.un395_half_pc_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__15937\,
            in1 => \N__21456\,
            in2 => \N__12464\,
            in3 => \N__27641\,
            lcout => \processor_zipi8.program_counter_i.un395_half_pcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIQQO068_7_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010100000000"
        )
    port map (
            in0 => \N__14236\,
            in1 => \N__15935\,
            in2 => \N__14261\,
            in3 => \N__14267\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_46_7\,
            ltout => \processor_zipi8.program_counter_i.carry_pc_46_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIT0QD69_8_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__15936\,
            in1 => \N__13049\,
            in2 => \N__13040\,
            in3 => \N__12874\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_52_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNI8JKGO_8_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__17775\,
            in1 => \N__17860\,
            in2 => \N__12943\,
            in3 => \N__21111\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNO_0_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__16889\,
            in1 => \N__12836\,
            in2 => \N__12860\,
            in3 => \N__17903\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.zero_flag_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__17400\,
            in1 => \N__17506\,
            in2 => \N__12863\,
            in3 => \N__18033\,
            lcout => \processor_zipi8.zero_flag\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33633\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.shadow_zero_flag_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12809\,
            lcout => \processor_zipi8.shadow_zero_flag\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33633\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_6_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34083\,
            in1 => \N__29371\,
            in2 => \N__29736\,
            in3 => \N__35861\,
            lcout => OPEN,
            ltout => \processor_zipi8.alu_result_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNO_1_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12851\,
            in1 => \N__12830\,
            in2 => \N__12839\,
            in3 => \N__13091\,
            lcout => \processor_zipi8.flags_i.zero_flag_3_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_5_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34081\,
            in1 => \N__29952\,
            in2 => \N__30492\,
            in3 => \N__35859\,
            lcout => \processor_zipi8.alu_result_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.shadow_carry_flag_1_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12824\,
            lcout => \processor_zipi8.stack_i.shadow_zero_value\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33633\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_3_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34082\,
            in1 => \N__37628\,
            in2 => \N__38174\,
            in3 => \N__35860\,
            lcout => \processor_zipi8.alu_result_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI0LOT3_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14658\,
            in2 => \_gnd_net_\,
            in3 => \N__14325\,
            lcout => \processor_zipi8.flags_i.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNICAJR_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__18029\,
            in1 => \N__17989\,
            in2 => \_gnd_net_\,
            in3 => \N__24112\,
            lcout => \processor_zipi8.flags_i.m49_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIJK644_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100001000"
        )
    port map (
            in0 => \N__14327\,
            in1 => \N__19042\,
            in2 => \N__16290\,
            in3 => \N__14660\,
            lcout => \processor_zipi8.flags_i.m82_1\,
            ltout => \processor_zipi8.flags_i.m82_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.stack_pointer_1_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__14560\,
            in1 => \N__17394\,
            in2 => \N__13085\,
            in3 => \N__16276\,
            lcout => \processor_zipi8.stack_pointer_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIJSPM4_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__16275\,
            in1 => \N__13082\,
            in2 => \N__17416\,
            in3 => \N__14559\,
            lcout => \processor_zipi8.zero_flag_RNIJSPM4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIALV04_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14659\,
            in1 => \N__16271\,
            in2 => \_gnd_net_\,
            in3 => \N__14326\,
            lcout => \processor_zipi8.flags_i.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI6N578_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__14486\,
            in1 => \N__14455\,
            in2 => \N__15167\,
            in3 => \N__13058\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.m61_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNID5QI8_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100101"
        )
    port map (
            in0 => \N__15165\,
            in1 => \N__17260\,
            in2 => \N__13052\,
            in3 => \N__16280\,
            lcout => \processor_zipi8.flags_i.i14_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI3VC94_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000110101"
        )
    port map (
            in0 => \N__14456\,
            in1 => \N__14661\,
            in2 => \N__16291\,
            in3 => \N__14487\,
            lcout => \processor_zipi8.flags_i.zero_flag_RNI3VCZ0Z94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__7_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34520\,
            in1 => \N__36661\,
            in2 => \N__33013\,
            in3 => \N__33316\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33642\,
            ce => \N__26167\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNITSK21_6_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__13130\,
            in1 => \N__31745\,
            in2 => \N__16445\,
            in3 => \N__30985\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIGUSR1_6_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__13262\,
            in1 => \N__31744\,
            in2 => \N__13133\,
            in3 => \N__16394\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIGUSR1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_6_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16441\,
            in1 => \N__13129\,
            in2 => \_gnd_net_\,
            in3 => \N__37468\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__6_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34303\,
            in1 => \N__36557\,
            in2 => \N__29365\,
            in3 => \N__29706\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33636\,
            ce => \N__18076\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_6_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16393\,
            in1 => \N__13261\,
            in2 => \_gnd_net_\,
            in3 => \N__37467\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIVUK21_7_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30986\,
            in1 => \N__16427\,
            in2 => \N__31751\,
            in3 => \N__13103\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIK2TR1_7_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__16541\,
            in2 => \N__13118\,
            in3 => \N__31749\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIK2TR1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__7_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34304\,
            in1 => \N__32978\,
            in2 => \N__33359\,
            in3 => \N__36558\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33636\,
            ce => \N__18076\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_6_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13210\,
            in1 => \N__37394\,
            in2 => \_gnd_net_\,
            in3 => \N__16483\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI70021_6_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__16484\,
            in1 => \N__31698\,
            in2 => \N__31014\,
            in3 => \N__13211\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNII1NP1_6_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__13430\,
            in1 => \N__31701\,
            in2 => \N__13190\,
            in3 => \N__13316\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNII1NP1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_6_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37395\,
            in1 => \N__13315\,
            in2 => \_gnd_net_\,
            in3 => \N__13429\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_6_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__13187\,
            in1 => \N__28649\,
            in2 => \N__13181\,
            in3 => \N__29012\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_6_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28650\,
            in1 => \N__13178\,
            in2 => \N__13169\,
            in3 => \N__13166\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_6_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__14753\,
            in1 => \N__25667\,
            in2 => \N__13157\,
            in3 => \N__25785\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_6_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25668\,
            in1 => \N__23828\,
            in2 => \N__13154\,
            in3 => \N__24611\,
            lcout => \processor_zipi8.sy_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34751\,
            in1 => \N__36553\,
            in2 => \N__32460\,
            in3 => \N__32026\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__36549\,
            in1 => \N__34756\,
            in2 => \N__39233\,
            in3 => \N__39592\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__2_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__38556\,
            in1 => \N__36554\,
            in2 => \N__34840\,
            in3 => \N__38730\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__3_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36550\,
            in1 => \N__34754\,
            in2 => \N__38184\,
            in3 => \N__37825\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__4_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34752\,
            in1 => \N__36555\,
            in2 => \N__35560\,
            in3 => \N__35156\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__5_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36551\,
            in1 => \N__34755\,
            in2 => \N__30499\,
            in3 => \N__29951\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__6_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34753\,
            in1 => \N__36556\,
            in2 => \N__29705\,
            in3 => \N__29315\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__7_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36552\,
            in1 => \N__33271\,
            in2 => \N__32995\,
            in3 => \N__34760\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33625\,
            ce => \N__14876\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34556\,
            in1 => \N__36596\,
            in2 => \N__32433\,
            in3 => \N__32025\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33616\,
            ce => \N__20288\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__2_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36593\,
            in1 => \N__34558\,
            in2 => \N__38802\,
            in3 => \N__38557\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33616\,
            ce => \N__20288\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__3_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__37774\,
            in1 => \N__38154\,
            in2 => \N__34764\,
            in3 => \N__36598\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33616\,
            ce => \N__20288\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__5_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36594\,
            in1 => \N__34559\,
            in2 => \N__30508\,
            in3 => \N__29950\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33616\,
            ce => \N__20288\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_5_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18296\,
            in1 => \N__18274\,
            in2 => \_gnd_net_\,
            in3 => \N__37484\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__6_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36595\,
            in1 => \N__34560\,
            in2 => \N__29770\,
            in3 => \N__29316\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33616\,
            ce => \N__20288\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__7_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34557\,
            in1 => \N__36597\,
            in2 => \N__33017\,
            in3 => \N__33319\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33616\,
            ce => \N__20288\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_7_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37485\,
            in1 => \N__16537\,
            in2 => \_gnd_net_\,
            in3 => \N__13243\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34742\,
            in1 => \N__36370\,
            in2 => \N__32432\,
            in3 => \N__32024\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__1_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36366\,
            in1 => \N__34745\,
            in2 => \N__39598\,
            in3 => \N__39224\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__2_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__38513\,
            in1 => \N__36371\,
            in2 => \N__34839\,
            in3 => \N__38729\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__3_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__36367\,
            in1 => \N__34747\,
            in2 => \N__37862\,
            in3 => \N__38147\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__4_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34743\,
            in1 => \N__36372\,
            in2 => \N__35211\,
            in3 => \N__35573\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__5_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36368\,
            in1 => \N__34746\,
            in2 => \N__30444\,
            in3 => \N__29894\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__6_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34744\,
            in1 => \N__29311\,
            in2 => \N__29769\,
            in3 => \N__36373\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__7_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__36369\,
            in1 => \N__33318\,
            in2 => \N__34841\,
            in3 => \N__32993\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33610\,
            ce => \N__14897\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34402\,
            in1 => \N__36201\,
            in2 => \N__32431\,
            in3 => \N__32023\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33607\,
            ce => \N__14863\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36197\,
            in1 => \N__39545\,
            in2 => \N__39228\,
            in3 => \N__34406\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33607\,
            ce => \N__14863\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__2_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34403\,
            in1 => \N__36202\,
            in2 => \N__38558\,
            in3 => \N__38725\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33607\,
            ce => \N__14863\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__3_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36198\,
            in1 => \N__34405\,
            in2 => \N__38185\,
            in3 => \N__37797\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33607\,
            ce => \N__14863\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_5_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14912\,
            in1 => \N__13289\,
            in2 => \_gnd_net_\,
            in3 => \N__36196\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202\,
            ltout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__5_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36199\,
            in1 => \N__30461\,
            in2 => \N__13283\,
            in3 => \N__34407\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33607\,
            ce => \N__14863\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__4_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34404\,
            in1 => \N__35155\,
            in2 => \N__35569\,
            in3 => \N__36203\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33607\,
            ce => \N__14863\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__6_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36200\,
            in1 => \N__29684\,
            in2 => \N__29366\,
            in3 => \N__34408\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33607\,
            ce => \N__14863\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_6_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__13351\,
            in1 => \N__19474\,
            in2 => \N__16633\,
            in3 => \N__19798\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_6_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13331\,
            in1 => \N__13376\,
            in2 => \N__13415\,
            in3 => \N__13412\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_6_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101111111"
        )
    port map (
            in0 => \N__19640\,
            in1 => \N__16630\,
            in2 => \N__13362\,
            in3 => \N__19587\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_1_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28652\,
            in1 => \_gnd_net_\,
            in2 => \N__21458\,
            in3 => \N__13405\,
            lcout => \processor_zipi8.port_id_6\,
            ltout => \processor_zipi8.port_id_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_6_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__16623\,
            in1 => \N__19586\,
            in2 => \N__13379\,
            in3 => \N__19206\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_6_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110111"
        )
    port map (
            in0 => \N__19205\,
            in1 => \N__13355\,
            in2 => \N__16634\,
            in3 => \N__24012\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIF3G21_6_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13520\,
            in1 => \N__21448\,
            in2 => \_gnd_net_\,
            in3 => \N__28651\,
            lcout => \processor_zipi8.pc_vector_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_6_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13529\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.state_machine_i.t_state_1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__17339\,
            in1 => \N__19005\,
            in2 => \N__13460\,
            in3 => \N__16289\,
            lcout => \processor_zipi8.t_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_2_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16868\,
            in2 => \_gnd_net_\,
            in3 => \N__17021\,
            lcout => \processor_zipi8.arith_logical_result_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m38_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__13486\,
            in1 => \N__13879\,
            in2 => \_gnd_net_\,
            in3 => \N__15144\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.N_125_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.state_machine_i.run_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13501\,
            in2 => \N__13511\,
            in3 => \N__17340\,
            lcout => \processor_zipi8.run\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.shadow_carry_flag_3_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13508\,
            lcout => \processor_zipi8.special_bit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.state_machine_i.internal_reset_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101110011"
        )
    port map (
            in0 => \N__13880\,
            in1 => \N__13500\,
            in2 => \N__15158\,
            in3 => \N__13487\,
            lcout => \processor_zipi8.internal_reset\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_2_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13466\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.state_machine_i.t_state_2_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__16288\,
            in1 => \N__13459\,
            in2 => \N__19041\,
            in3 => \N__17341\,
            lcout => \processor_zipi8.state_machine_i.bram_enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_11_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13436\,
            lcout => \processor_zipi8.return_vector_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m36_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111011111"
        )
    port map (
            in0 => \N__17255\,
            in1 => \N__19000\,
            in2 => \N__15113\,
            in3 => \N__16287\,
            lcout => \processor_zipi8.flags_i.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.stack_pointer_4_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__19001\,
            in1 => \N__15827\,
            in2 => \N__17379\,
            in3 => \N__15803\,
            lcout => \processor_zipi8.stack_pointer_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_7_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13871\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_1_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13859\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINQ3G8_5_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__13847\,
            in1 => \N__23663\,
            in2 => \N__18263\,
            in3 => \N__27316\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5QUHH_5_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22790\,
            in2 => \N__13835\,
            in3 => \N__22232\,
            lcout => \processor_zipi8.sx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_4_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101100110011001"
        )
    port map (
            in0 => \N__15332\,
            in1 => \N__13535\,
            in2 => \N__15954\,
            in3 => \N__21245\,
            lcout => address_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33627\,
            ce => \N__15762\,
            sr => \N__17444\
        );

    \processor_zipi8.program_counter_i.pc_esr_6_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101001010101"
        )
    port map (
            in0 => \N__14303\,
            in1 => \N__15933\,
            in2 => \N__14297\,
            in3 => \N__14276\,
            lcout => address_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33627\,
            ce => \N__15762\,
            sr => \N__17444\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIJE19O_4_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__17881\,
            in1 => \N__16948\,
            in2 => \N__13586\,
            in3 => \N__17799\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_4\,
            ltout => \processor_zipi8.program_counter_i.half_pc_0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIBG8G55_4_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100000000"
        )
    port map (
            in0 => \N__21244\,
            in1 => \N__15926\,
            in2 => \N__14309\,
            in3 => \N__15331\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_28_4\,
            ltout => \processor_zipi8.program_counter_i.carry_pc_28_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIOGNL56_5_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__15927\,
            in1 => \N__14059\,
            in2 => \N__14306\,
            in3 => \N__14074\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_34_5\,
            ltout => \processor_zipi8.program_counter_i.carry_pc_34_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNI8K7R57_6_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__14293\,
            in1 => \N__15928\,
            in2 => \N__14279\,
            in3 => \N__14275\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_40_6\,
            ltout => \processor_zipi8.program_counter_i.carry_pc_40_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_7_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000001111"
        )
    port map (
            in0 => \N__15934\,
            in1 => \N__14260\,
            in2 => \N__14240\,
            in3 => \N__14237\,
            lcout => address_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33627\,
            ce => \N__15762\,
            sr => \N__17444\
        );

    \processor_zipi8.program_counter_i.pc_esr_5_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101011010101"
        )
    port map (
            in0 => \N__14075\,
            in1 => \N__15932\,
            in2 => \N__14063\,
            in3 => \N__14048\,
            lcout => address_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33627\,
            ce => \N__15762\,
            sr => \N__17444\
        );

    \processor_zipi8.program_counter_i.un3_half_pc_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17857\,
            in2 => \_gnd_net_\,
            in3 => \N__17771\,
            lcout => \processor_zipi8.program_counter_i.un3_half_pcZ0\,
            ltout => \processor_zipi8.program_counter_i.un3_half_pcZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNO_1_11_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__13892\,
            in1 => \N__21432\,
            in2 => \N__13883\,
            in3 => \N__27442\,
            lcout => \processor_zipi8.program_counter_i.un431_half_pc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNIKAV8O_2_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__15227\,
            in1 => \N__17773\,
            in2 => \N__25540\,
            in3 => \N__17859\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNO_0_11_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__20051\,
            in1 => \N__14398\,
            in2 => \N__17871\,
            in3 => \N__17774\,
            lcout => OPEN,
            ltout => \processor_zipi8.program_counter_i.half_pc_0_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_11_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101011001111"
        )
    port map (
            in0 => \N__14417\,
            in1 => \N__14411\,
            in2 => \N__14405\,
            in3 => \N__14353\,
            lcout => \processor_zipi8.address_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33635\,
            ce => \N__15767\,
            sr => \N__17425\
        );

    \processor_zipi8.program_counter_i.pc_RNI70TDO_0_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011101110"
        )
    port map (
            in0 => \N__15449\,
            in1 => \N__17772\,
            in2 => \N__23012\,
            in3 => \N__17858\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNI2ASQ6A_9_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010100000000"
        )
    port map (
            in0 => \N__14387\,
            in1 => \N__15938\,
            in2 => \N__14381\,
            in3 => \N__14365\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_58_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIJJ175_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__21179\,
            in1 => \N__14423\,
            in2 => \N__18908\,
            in3 => \N__14432\,
            lcout => \processor_zipi8.pc_mode_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIOK4K1_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011100010010"
        )
    port map (
            in0 => \N__19932\,
            in1 => \N__14567\,
            in2 => \N__14342\,
            in3 => \N__21443\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.N_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI7M013_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14315\,
            in2 => \N__14333\,
            in3 => \N__24308\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.N_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIK0IP3_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010001"
        )
    port map (
            in0 => \N__14569\,
            in1 => \N__18874\,
            in2 => \N__14330\,
            in3 => \N__21180\,
            lcout => \processor_zipi8.flags_i.N_123_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m44_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111110101010"
        )
    port map (
            in0 => \N__21442\,
            in1 => \N__19931\,
            in2 => \N__14577\,
            in3 => \N__24172\,
            lcout => \processor_zipi8.flags_i.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m91_am_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001100110"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__14568\,
            in2 => \N__19958\,
            in3 => \N__21444\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.m91_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNINARM2_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__14714\,
            in1 => \_gnd_net_\,
            in2 => \N__14441\,
            in3 => \N__24309\,
            lcout => \processor_zipi8.flags_i.N_1239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m33_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14491\,
            in1 => \N__16270\,
            in2 => \N__14578\,
            in3 => \N__14657\,
            lcout => \processor_zipi8.flags_i.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNICAJR_0_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__18023\,
            in1 => \N__24094\,
            in2 => \_gnd_net_\,
            in3 => \N__17984\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.m25_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNID1UF1_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21437\,
            in2 => \N__14438\,
            in3 => \N__19901\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.N_26_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI04EE2_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010001"
        )
    port map (
            in0 => \N__21438\,
            in1 => \N__24096\,
            in2 => \N__14435\,
            in3 => \N__24293\,
            lcout => \processor_zipi8.flags_i.N_27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIULO51_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100101011101"
        )
    port map (
            in0 => \N__24095\,
            in1 => \N__24291\,
            in2 => \N__17993\,
            in3 => \N__18024\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.m20_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIHO842_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111110100"
        )
    port map (
            in0 => \N__19902\,
            in1 => \N__21439\,
            in2 => \N__14426\,
            in3 => \N__24292\,
            lcout => \processor_zipi8.flags_i.N_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m87_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14553\,
            in2 => \_gnd_net_\,
            in3 => \N__19903\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.N_1235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI89V91_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011010010"
        )
    port map (
            in0 => \N__18025\,
            in1 => \N__24097\,
            in2 => \N__14717\,
            in3 => \N__17988\,
            lcout => \processor_zipi8.flags_i.zero_flag_RNI89VZ0Z91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI4LCF3_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010001"
        )
    port map (
            in0 => \N__14554\,
            in1 => \N__18913\,
            in2 => \N__14708\,
            in3 => \N__21211\,
            lcout => \processor_zipi8.flags_i.N_124_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI281Q3_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011000000110"
        )
    port map (
            in0 => \N__14555\,
            in1 => \N__16278\,
            in2 => \N__19069\,
            in3 => \N__14699\,
            lcout => \processor_zipi8.flags_i.N_1241\,
            ltout => \processor_zipi8.flags_i.N_1241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIDS654_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__17402\,
            in1 => \_gnd_net_\,
            in2 => \N__14693\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.zero_flag_RNIDS654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.stack_pointer_2_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__19057\,
            in1 => \N__17405\,
            in2 => \N__14624\,
            in3 => \N__14612\,
            lcout => \processor_zipi8.stack_pointer_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m75_am_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__16279\,
            in1 => \N__14662\,
            in2 => \N__14573\,
            in3 => \N__14485\,
            lcout => \processor_zipi8.flags_i.m75_amZ0\,
            ltout => \processor_zipi8.flags_i.m75_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI5GK75_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__19056\,
            in1 => \N__17403\,
            in2 => \N__14615\,
            in3 => \N__14611\,
            lcout => \processor_zipi8.zero_flag_RNI5GK75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.stack_pointer_0_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14588\,
            lcout => \processor_zipi8.stack_pointer_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNI51D94_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001000111"
        )
    port map (
            in0 => \N__14484\,
            in1 => \N__16277\,
            in2 => \N__17259\,
            in3 => \N__14454\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.m68_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIAKL05_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010110001"
        )
    port map (
            in0 => \N__19009\,
            in1 => \N__17251\,
            in2 => \N__14759\,
            in3 => \N__15102\,
            lcout => \processor_zipi8.flags_i.N_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__6_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34128\,
            in1 => \N__36503\,
            in2 => \N__29329\,
            in3 => \N__29677\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33654\,
            ce => \N__23563\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__7_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36502\,
            in1 => \N__33311\,
            in2 => \N__33009\,
            in3 => \N__34129\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33654\,
            ce => \N__23563\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__6_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34305\,
            in1 => \N__29201\,
            in2 => \N__36626\,
            in3 => \N__29676\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33648\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_6_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16360\,
            in1 => \N__22376\,
            in2 => \_gnd_net_\,
            in3 => \N__37384\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_6_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__14831\,
            in1 => \N__14735\,
            in2 => \N__14756\,
            in3 => \N__28620\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_6_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16111\,
            in1 => \N__16093\,
            in2 => \_gnd_net_\,
            in3 => \N__37381\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_6_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37382\,
            in1 => \N__23809\,
            in2 => \_gnd_net_\,
            in3 => \N__16123\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_6_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__28619\,
            in1 => \N__14744\,
            in2 => \N__14738\,
            in3 => \N__29002\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_6_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14921\,
            in1 => \N__14729\,
            in2 => \_gnd_net_\,
            in3 => \N__36034\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268\,
            ltout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__6_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34127\,
            in1 => \N__29691\,
            in2 => \N__14834\,
            in3 => \N__36455\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33644\,
            ce => \N__25335\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_6_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37383\,
            in1 => \_gnd_net_\,
            in2 => \N__23462\,
            in3 => \N__16378\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_0_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14824\,
            in1 => \N__37078\,
            in2 => \_gnd_net_\,
            in3 => \N__14809\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIRJV11_0_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__16510\,
            in1 => \N__30922\,
            in2 => \N__31742\,
            in3 => \N__14792\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIQ8MP1_0_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__14825\,
            in1 => \N__14810\,
            in2 => \N__14795\,
            in3 => \N__31717\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIQ8MP1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_0_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37081\,
            in1 => \_gnd_net_\,
            in2 => \N__16511\,
            in3 => \N__14791\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__28617\,
            in1 => \N__28978\,
            in2 => \N__14777\,
            in3 => \N__14774\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_0_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__14765\,
            in1 => \N__14882\,
            in2 => \N__14768\,
            in3 => \N__28618\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_0_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18139\,
            in2 => \N__18121\,
            in3 => \N__37079\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_0_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37080\,
            in1 => \N__20387\,
            in2 => \_gnd_net_\,
            in3 => \N__20368\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe13_0_a2_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20856\,
            in1 => \N__22246\,
            in2 => \N__27461\,
            in3 => \N__20540\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe16_0_a2_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27445\,
            in1 => \N__23153\,
            in2 => \N__22284\,
            in3 => \N__20854\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20855\,
            in1 => \N__22245\,
            in2 => \N__20326\,
            in3 => \N__27447\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe8_0_a2_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27449\,
            in1 => \N__23159\,
            in2 => \N__22287\,
            in3 => \N__20857\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe10_0_a2_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20657\,
            in1 => \N__22247\,
            in2 => \N__23163\,
            in3 => \N__27448\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe18_0_a2_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27443\,
            in1 => \N__23154\,
            in2 => \N__22286\,
            in3 => \N__20658\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20659\,
            in1 => \N__22241\,
            in2 => \N__23164\,
            in3 => \N__27446\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe2_0_a2_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27444\,
            in1 => \N__23158\,
            in2 => \N__22285\,
            in3 => \N__20660\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe11_0_a2_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22138\,
            in1 => \N__20627\,
            in2 => \N__20324\,
            in3 => \N__27455\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe23_0_a2_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27451\,
            in1 => \N__20539\,
            in2 => \N__20646\,
            in3 => \N__22135\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe17_0_a2_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22134\,
            in1 => \N__20842\,
            in2 => \N__20325\,
            in3 => \N__27453\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe27_0_a2_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27452\,
            in1 => \N__20316\,
            in2 => \N__20647\,
            in3 => \N__22136\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe15_0_a2_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22137\,
            in1 => \N__20628\,
            in2 => \N__20543\,
            in3 => \N__27454\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe9_0_a2_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__27456\,
            in1 => \N__22139\,
            in2 => \N__20858\,
            in3 => \N__20317\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_0_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27631\,
            in2 => \_gnd_net_\,
            in3 => \N__30984\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212\,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe1_0_a2_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__27450\,
            in1 => \N__20841\,
            in2 => \N__14885\,
            in3 => \N__22133\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__21702\,
            in1 => \N__14932\,
            in2 => \_gnd_net_\,
            in3 => \N__17129\,
            lcout => \processor_zipi8.shift_rotate_result_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_2_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17128\,
            in1 => \N__20052\,
            in2 => \_gnd_net_\,
            in3 => \N__21701\,
            lcout => \processor_zipi8.shift_rotate_result_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_4_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17127\,
            in2 => \N__20057\,
            in3 => \N__18801\,
            lcout => \processor_zipi8.shift_rotate_result_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_6_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17125\,
            in1 => \N__16694\,
            in2 => \_gnd_net_\,
            in3 => \N__18802\,
            lcout => \processor_zipi8.shift_rotate_result_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_7_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__17124\,
            in1 => \N__16615\,
            in2 => \_gnd_net_\,
            in3 => \N__14933\,
            lcout => \processor_zipi8.shift_rotate_result_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_5_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17122\,
            in2 => \N__16631\,
            in3 => \N__21856\,
            lcout => \processor_zipi8.shift_rotate_result_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_3_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21855\,
            in1 => \N__17126\,
            in2 => \_gnd_net_\,
            in3 => \N__22044\,
            lcout => \processor_zipi8.shift_rotate_result_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22045\,
            in1 => \N__17123\,
            in2 => \_gnd_net_\,
            in3 => \N__21106\,
            lcout => \processor_zipi8.shift_rotate_result_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33612\,
            ce => 'H',
            sr => \N__25796\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_5_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14969\,
            in1 => \N__21441\,
            in2 => \_gnd_net_\,
            in3 => \N__25541\,
            lcout => \processor_zipi8.port_id_2\,
            ltout => \processor_zipi8.port_id_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_2_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101011111"
        )
    port map (
            in0 => \N__19577\,
            in1 => \N__19618\,
            in2 => \N__14900\,
            in3 => \N__22040\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__22041\,
            in1 => \N__19578\,
            in2 => \N__15045\,
            in3 => \N__19180\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_2_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__15034\,
            in1 => \N__23999\,
            in2 => \N__19202\,
            in3 => \N__22042\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_2_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111111111111"
        )
    port map (
            in0 => \N__22039\,
            in1 => \N__19794\,
            in2 => \N__19487\,
            in3 => \N__15035\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15011\,
            in1 => \N__15005\,
            in2 => \N__14999\,
            in3 => \N__14996\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI9VF21_2_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14990\,
            in1 => \N__14968\,
            in2 => \_gnd_net_\,
            in3 => \N__21440\,
            lcout => \processor_zipi8.pc_vector_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_RNO_5_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110100101"
        )
    port map (
            in0 => \N__32324\,
            in1 => \N__21227\,
            in2 => \N__39546\,
            in3 => \N__17990\,
            lcout => \processor_zipi8.flags_i.parity_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_3_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001011111101"
        )
    port map (
            in0 => \N__15350\,
            in1 => \N__15371\,
            in2 => \N__15980\,
            in3 => \N__15869\,
            lcout => address_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33630\,
            ce => \N__15758\,
            sr => \N__17390\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110111111101"
        )
    port map (
            in0 => \N__17991\,
            in1 => \N__21516\,
            in2 => \N__14975\,
            in3 => \N__17002\,
            lcout => OPEN,
            ltout => \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_1_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__21517\,
            in1 => \N__16702\,
            in2 => \N__14978\,
            in3 => \N__14973\,
            lcout => OPEN,
            ltout => \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__14974\,
            in1 => \N__21518\,
            in2 => \N__14936\,
            in3 => \N__21090\,
            lcout => \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.register_bank_control_i.bank_RNO_1_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__16049\,
            in1 => \N__17543\,
            in2 => \N__19059\,
            in3 => \N__16718\,
            lcout => \processor_zipi8.register_bank_control_i.un1_bank_value\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_2_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000110011"
        )
    port map (
            in0 => \N__15370\,
            in1 => \N__15976\,
            in2 => \_gnd_net_\,
            in3 => \N__15349\,
            lcout => address_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33630\,
            ce => \N__15758\,
            sr => \N__17390\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5LPHH_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22132\,
            in1 => \N__24779\,
            in2 => \_gnd_net_\,
            in3 => \N__20555\,
            lcout => \processor_zipi8.sx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m57_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__17230\,
            in1 => \N__15157\,
            in2 => \_gnd_net_\,
            in3 => \N__15109\,
            lcout => \processor_zipi8.flags_i.i14_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_RNO_0_0_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101100000000"
        )
    port map (
            in0 => \N__16013\,
            in1 => \N__15956\,
            in2 => \N__15062\,
            in3 => \N__15842\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_7_0_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21401\,
            in1 => \N__17000\,
            in2 => \_gnd_net_\,
            in3 => \N__23005\,
            lcout => \processor_zipi8.port_id_0\,
            ltout => \processor_zipi8.port_id_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101111111"
        )
    port map (
            in0 => \N__19457\,
            in1 => \N__19783\,
            in2 => \N__15083\,
            in3 => \N__21083\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_1_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17030\,
            in2 => \_gnd_net_\,
            in3 => \N__19283\,
            lcout => \processor_zipi8.arith_logical_result_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_0_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15080\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI6TF21_0_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21402\,
            in1 => \N__15068\,
            in2 => \_gnd_net_\,
            in3 => \N__17001\,
            lcout => \processor_zipi8.pc_vector_0\,
            ltout => \processor_zipi8.pc_vector_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_RNIUJNL41_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100000000"
        )
    port map (
            in0 => \N__16012\,
            in1 => \N__15955\,
            in2 => \N__15845\,
            in3 => \N__15841\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNIC4FP9_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000101"
        )
    port map (
            in0 => \N__17414\,
            in1 => \N__19066\,
            in2 => \N__15826\,
            in3 => \N__15802\,
            lcout => \processor_zipi8.zero_flag_RNIC4FP9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_ctle_11_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17412\,
            in2 => \_gnd_net_\,
            in3 => \N__19065\,
            lcout => \processor_zipi8.program_counter_i.t_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_RNI72UDO_1_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010111001111"
        )
    port map (
            in0 => \N__17850\,
            in1 => \N__17798\,
            in2 => \N__15611\,
            in3 => \N__23198\,
            lcout => OPEN,
            ltout => \processor_zipi8.program_counter_i.half_pc_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_RNINDAA01_1_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21482\,
            in2 => \N__15722\,
            in3 => \N__15957\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_1\,
            ltout => \processor_zipi8.program_counter_i.half_pc_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_1_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__15348\,
            in1 => \N__15602\,
            in2 => \N__15719\,
            in3 => \N__19068\,
            lcout => address_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33643\,
            ce => 'H',
            sr => \N__17415\
        );

    \processor_zipi8.program_counter_i.pc_0_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__19067\,
            in1 => \N__15548\,
            in2 => \_gnd_net_\,
            in3 => \N__15441\,
            lcout => address_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33643\,
            ce => 'H',
            sr => \N__17415\
        );

    \processor_zipi8.flags_i.zero_flag_RNIL8RB5_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__17413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17281\,
            lcout => \processor_zipi8.zero_flag_RNIL8RB5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNI3JQA54_3_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__15970\,
            in1 => \N__15865\,
            in2 => \N__15369\,
            in3 => \N__15347\,
            lcout => \processor_zipi8.program_counter_i.carry_pc_22_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__24153\,
            in1 => \N__16730\,
            in2 => \N__18883\,
            in3 => \N__24276\,
            lcout => \processor_zipi8.pc_mode_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNI6NB501_2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__15998\,
            in1 => \N__15958\,
            in2 => \_gnd_net_\,
            in3 => \N__15989\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNI8QC501_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__15959\,
            in1 => \N__17054\,
            in2 => \_gnd_net_\,
            in3 => \N__17573\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.arith_logical_sel_1_1_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__24275\,
            in1 => \N__19944\,
            in2 => \_gnd_net_\,
            in3 => \N__24154\,
            lcout => \processor_zipi8.arith_logical_sel_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m101_e_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__24155\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24277\,
            lcout => \processor_zipi8.un16_alu_mux_sel_value\,
            ltout => \processor_zipi8.un16_alu_mux_sel_value_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.register_bank_control_i.sx_addr_4_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__16133\,
            in1 => \_gnd_net_\,
            in2 => \N__15854\,
            in3 => \N__25609\,
            lcout => \processor_zipi8.sx_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_4_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__21216\,
            in1 => \N__24161\,
            in2 => \N__18884\,
            in3 => \N__24278\,
            lcout => \processor_zipi8.decode4_strobes_enables_i.un23_flag_enable_type\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_pc_statck_i.returni_type_o_2_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21215\,
            in2 => \_gnd_net_\,
            in3 => \N__19945\,
            lcout => \processor_zipi8.returni_type_o_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_3_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__21224\,
            in1 => \N__19937\,
            in2 => \N__18931\,
            in3 => \N__15851\,
            lcout => OPEN,
            ltout => \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_1_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__19938\,
            in1 => \N__18921\,
            in2 => \N__16076\,
            in3 => \N__24289\,
            lcout => \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_2_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16073\,
            in1 => \N__16064\,
            in2 => \_gnd_net_\,
            in3 => \N__35731\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.register_bank_control_i.bank_RNO_4_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19936\,
            in1 => \N__21223\,
            in2 => \N__21457\,
            in3 => \N__24288\,
            lcout => OPEN,
            ltout => \processor_zipi8.register_bank_control_i.un31_regbank_type_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.register_bank_control_i.bank_RNO_3_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18914\,
            in2 => \N__16052\,
            in3 => \N__24170\,
            lcout => \processor_zipi8.register_bank_control_i.un31_regbank_type\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.spm_enable_RNO_0_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19939\,
            in1 => \N__21225\,
            in2 => \N__18930\,
            in3 => \N__19060\,
            lcout => \processor_zipi8.decode4_strobes_enables_i.spm_enable_value_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_0_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16040\,
            in1 => \N__35730\,
            in2 => \_gnd_net_\,
            in3 => \N__16031\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.alu_mux_sel_1_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__24171\,
            in1 => \_gnd_net_\,
            in2 => \N__19959\,
            in3 => \N__24290\,
            lcout => \processor_zipi8.alu_mux_sel_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__16304\,
            in1 => \N__17924\,
            in2 => \N__18929\,
            in3 => \N__24331\,
            lcout => OPEN,
            ltout => \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16016\,
            in3 => \N__16298\,
            lcout => \processor_zipi8.pc_mode_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_pc_statck_i.un3_pc_mode_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__21416\,
            in1 => \N__24327\,
            in2 => \N__24169\,
            in3 => \N__21181\,
            lcout => \processor_zipi8.decode4_pc_statck_i.un3_pc_modeZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m16_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__24147\,
            in1 => \N__21417\,
            in2 => \N__24340\,
            in3 => \N__19946\,
            lcout => \processor_zipi8.N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.m104_2_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__21182\,
            in1 => \N__18912\,
            in2 => \N__16292\,
            in3 => \N__19947\,
            lcout => \processor_zipi8.flags_i.m104Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__7_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36688\,
            in1 => \N__34571\,
            in2 => \N__33342\,
            in3 => \N__33016\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33668\,
            ce => \N__24917\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__6_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34130\,
            in1 => \N__36484\,
            in2 => \N__29367\,
            in3 => \N__29675\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33662\,
            ce => \N__20141\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__7_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34569\,
            in1 => \N__33309\,
            in2 => \N__33014\,
            in3 => \N__36501\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33662\,
            ce => \N__20141\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__4_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34306\,
            in1 => \N__35193\,
            in2 => \N__36848\,
            in3 => \N__35427\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33655\,
            ce => \N__32674\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNINVTE1_6_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__16124\,
            in1 => \N__31590\,
            in2 => \N__23813\,
            in3 => \N__30932\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI44F42_6_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31591\,
            in1 => \N__16112\,
            in2 => \N__16100\,
            in3 => \N__16097\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI44F42_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMVAG4_6_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__27386\,
            in1 => \N__16343\,
            in2 => \N__16079\,
            in3 => \N__27640\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIVVE01_6_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30931\,
            in1 => \N__23461\,
            in2 => \N__31695\,
            in3 => \N__16379\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIK4HN1_6_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__22375\,
            in1 => \N__16361\,
            in2 => \N__16346\,
            in3 => \N__31589\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIK4HN1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7B4G8_6_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__16337\,
            in1 => \N__16328\,
            in2 => \N__16322\,
            in3 => \N__27387\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7B4G8_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5RVHH_6_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22415\,
            in2 => \N__16307\,
            in3 => \N__22234\,
            lcout => \processor_zipi8.sx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__36705\,
            in1 => \N__33951\,
            in2 => \N__32098\,
            in3 => \N__32240\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__33947\,
            in1 => \N__36709\,
            in2 => \N__39262\,
            in3 => \N__39591\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__2_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36706\,
            in1 => \N__33952\,
            in2 => \N__38881\,
            in3 => \N__38462\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__3_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__33948\,
            in1 => \N__36710\,
            in2 => \N__37824\,
            in3 => \N__38098\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__4_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__36707\,
            in1 => \N__33954\,
            in2 => \N__35191\,
            in3 => \N__35549\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__5_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__33949\,
            in1 => \N__36711\,
            in2 => \N__30463\,
            in3 => \N__30076\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__6_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36708\,
            in1 => \N__33953\,
            in2 => \N__29704\,
            in3 => \N__29357\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__7_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__33950\,
            in1 => \N__36712\,
            in2 => \N__32994\,
            in3 => \N__33256\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33645\,
            ce => \N__16409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34499\,
            in1 => \N__32380\,
            in2 => \N__32097\,
            in3 => \N__36814\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__36807\,
            in1 => \N__39247\,
            in2 => \N__39593\,
            in3 => \N__34505\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34500\,
            in1 => \N__36811\,
            in2 => \N__38532\,
            in3 => \N__38886\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__3_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36808\,
            in1 => \N__34503\,
            in2 => \N__38158\,
            in3 => \N__37701\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34501\,
            in1 => \N__36812\,
            in2 => \N__35192\,
            in3 => \N__35426\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__5_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36809\,
            in1 => \N__30386\,
            in2 => \N__30137\,
            in3 => \N__34506\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__6_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34502\,
            in1 => \N__36813\,
            in2 => \N__29301\,
            in3 => \N__29554\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__7_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36810\,
            in1 => \N__33266\,
            in2 => \N__33012\,
            in3 => \N__34504\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33638\,
            ce => \N__16523\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34507\,
            in1 => \N__32244\,
            in2 => \N__32099\,
            in3 => \N__36699\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__1_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36692\,
            in1 => \N__34511\,
            in2 => \N__39597\,
            in3 => \N__39094\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__2_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34508\,
            in1 => \N__36698\,
            in2 => \N__38540\,
            in3 => \N__38851\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__3_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36693\,
            in1 => \N__38099\,
            in2 => \N__37853\,
            in3 => \N__34512\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__4_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34509\,
            in1 => \N__36696\,
            in2 => \N__35218\,
            in3 => \N__35511\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__5_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36694\,
            in1 => \N__30394\,
            in2 => \N__30044\,
            in3 => \N__34513\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__6_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34510\,
            in1 => \N__36697\,
            in2 => \N__29364\,
            in3 => \N__29553\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__7_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36695\,
            in1 => \N__33174\,
            in2 => \N__33029\,
            in3 => \N__34514\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33631\,
            ce => \N__16454\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__0_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34516\,
            in1 => \N__36413\,
            in2 => \N__32299\,
            in3 => \N__31988\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33621\,
            ce => \N__18083\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__1_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36410\,
            in1 => \N__34518\,
            in2 => \N__39594\,
            in3 => \N__39052\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33621\,
            ce => \N__18083\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__2_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__38545\,
            in1 => \N__36414\,
            in2 => \N__38880\,
            in3 => \N__34515\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33621\,
            ce => \N__18083\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__36411\,
            in1 => \N__38123\,
            in2 => \N__34700\,
            in3 => \N__37801\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33621\,
            ce => \N__18083\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__4_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__34517\,
            in1 => \N__35363\,
            in2 => \N__36607\,
            in3 => \N__35006\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33621\,
            ce => \N__18083\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__5_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36412\,
            in1 => \N__34519\,
            in2 => \N__30462\,
            in3 => \N__30057\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33621\,
            ce => \N__18083\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_3_0_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16949\,
            in1 => \N__21445\,
            in2 => \_gnd_net_\,
            in3 => \N__37486\,
            lcout => \processor_zipi8.port_id_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.arith_carry_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__19796\,
            in1 => \N__16553\,
            in2 => \N__16706\,
            in3 => \N__16562\,
            lcout => \processor_zipi8.flags_i.arith_carryZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical6_process_carry_arith_logical_40_6_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__16798\,
            in1 => \N__19795\,
            in2 => \N__16619\,
            in3 => \N__19330\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6\,
            ltout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_7_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16556\,
            in3 => \N__16552\,
            lcout => \processor_zipi8.arith_logical_result_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_6_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__16799\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19331\,
            lcout => \processor_zipi8.arith_logical_result_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_RNO_3_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111110111"
        )
    port map (
            in0 => \N__16769\,
            in1 => \N__16910\,
            in2 => \N__19964\,
            in3 => \N__16756\,
            lcout => OPEN,
            ltout => \processor_zipi8.flags_i.carry_flag_value_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_RNO_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000000000"
        )
    port map (
            in0 => \N__16712\,
            in1 => \N__16775\,
            in2 => \N__16784\,
            in3 => \N__16736\,
            lcout => \processor_zipi8.flags_i.carry_flag_value_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_RNO_1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29499\,
            in1 => \N__19304\,
            in2 => \N__33147\,
            in3 => \N__16781\,
            lcout => \processor_zipi8.flags_i.carry_flag_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_RNO_2_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000111111"
        )
    port map (
            in0 => \N__16768\,
            in1 => \N__16879\,
            in2 => \N__16757\,
            in3 => \N__23986\,
            lcout => \processor_zipi8.flags_i.carry_flag_value_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un52_half_arith_logical_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__19779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19186\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21399\,
            in2 => \_gnd_net_\,
            in3 => \N__19949\,
            lcout => \processor_zipi8.decode4_pc_statck_i.N_22_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.register_bank_control_i.bank_RNO_2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21400\,
            in1 => \N__24323\,
            in2 => \N__18932\,
            in3 => \N__24163\,
            lcout => \processor_zipi8.register_bank_control_i.un17_regbank_type_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_RNO_4_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__24164\,
            in1 => \_gnd_net_\,
            in2 => \N__24338\,
            in3 => \N__19951\,
            lcout => \processor_zipi8.flags_i.un17_carry_flag_value_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.alu_mux_sel_value_1_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__19950\,
            in1 => \N__24319\,
            in2 => \_gnd_net_\,
            in3 => \N__24162\,
            lcout => \processor_zipi8.alu_mux_sel_value_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_1_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__24165\,
            in1 => \_gnd_net_\,
            in2 => \N__24339\,
            in3 => \N__17542\,
            lcout => \processor_zipi8.decode4_strobes_enables_i.un8_register_enable_type\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical2_process_carry_arith_logical_16_2_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__19780\,
            in1 => \N__16861\,
            in2 => \N__22043\,
            in3 => \N__17014\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2\,
            ltout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical3_process_carry_arith_logical_22_3_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20050\,
            in1 => \N__19102\,
            in2 => \N__16850\,
            in3 => \N__19781\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_22_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_21_tz_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__19467\,
            in1 => \N__19187\,
            in2 => \_gnd_net_\,
            in3 => \N__21685\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.N_773_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110111111111"
        )
    port map (
            in0 => \N__19188\,
            in1 => \N__21078\,
            in2 => \N__19778\,
            in3 => \N__16821\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__21079\,
            in1 => \N__16823\,
            in2 => \N__16847\,
            in3 => \N__23988\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_0_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000001110000"
        )
    port map (
            in0 => \N__19557\,
            in1 => \N__21080\,
            in2 => \N__16844\,
            in3 => \N__16822\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un36_half_arith_logical_1_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16824\,
            in2 => \_gnd_net_\,
            in3 => \N__19189\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__19294\,
            in1 => \N__21081\,
            in2 => \N__17048\,
            in3 => \N__17039\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0\,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical0_process_carry_arith_logical_4_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110100011"
        )
    port map (
            in0 => \N__21082\,
            in1 => \N__17563\,
            in2 => \N__17033\,
            in3 => \N__19743\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0\,
            ltout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical1_process_carry_arith_logical_10_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__21686\,
            in1 => \N__19784\,
            in2 => \N__17024\,
            in3 => \N__19279\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.register_bank_control_i.bank_RNO_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__24314\,
            in1 => \N__16916\,
            in2 => \_gnd_net_\,
            in3 => \N__17003\,
            lcout => OPEN,
            ltout => \processor_zipi8.register_bank_control_i.bank_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.register_bank_control_i.bank_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000101110"
        )
    port map (
            in0 => \N__25605\,
            in1 => \N__16964\,
            in2 => \N__16952\,
            in3 => \N__17442\,
            lcout => \processor_zipi8.bank\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_4_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__19343\,
            in1 => \N__19970\,
            in2 => \N__24590\,
            in3 => \N__25604\,
            lcout => \processor_zipi8.sy_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.shadow_carry_flag_2_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16931\,
            lcout => \processor_zipi8.shadow_bank\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.calc_arith_logical_sel_process_un4_arith_logical_sel_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16903\,
            in2 => \_gnd_net_\,
            in3 => \N__19948\,
            lcout => \processor_zipi8.un4_arith_logical_sel\,
            ltout => \processor_zipi8.un4_arith_logical_sel_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.arith_carry_in_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__21214\,
            in1 => \N__23976\,
            in2 => \N__16892\,
            in3 => \N__17959\,
            lcout => \processor_zipi8.arith_carry_in_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000110010"
        )
    port map (
            in0 => \N__17960\,
            in1 => \N__17443\,
            in2 => \N__17507\,
            in3 => \N__17453\,
            lcout => \processor_zipi8.carry_flag\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.stack_i.stack_pointer_3_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17441\,
            in2 => \_gnd_net_\,
            in3 => \N__17285\,
            lcout => \processor_zipi8.stack_pointer_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_3_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001111111111"
        )
    port map (
            in0 => \N__19631\,
            in1 => \N__19551\,
            in2 => \N__20046\,
            in3 => \N__17156\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__17135\,
            in1 => \N__17201\,
            in2 => \N__17204\,
            in3 => \N__17192\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_3_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__19563\,
            in1 => \N__17155\,
            in2 => \N__20045\,
            in3 => \N__19153\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_4_0_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17101\,
            in1 => \N__21356\,
            in2 => \_gnd_net_\,
            in3 => \N__19652\,
            lcout => \processor_zipi8.port_id_3\,
            ltout => \processor_zipi8.port_id_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_3_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101111111"
        )
    port map (
            in0 => \N__19473\,
            in1 => \N__20014\,
            in2 => \N__17195\,
            in3 => \N__19739\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_3_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__19152\,
            in1 => \N__20024\,
            in2 => \N__17166\,
            in3 => \N__23985\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIA0G21_3_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21355\,
            in1 => \N__23633\,
            in2 => \_gnd_net_\,
            in3 => \N__17100\,
            lcout => \processor_zipi8.pc_vector_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.program_counter_i.pc_esr_RNILC09O_3_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010111001111"
        )
    port map (
            in0 => \N__17849\,
            in1 => \N__17804\,
            in2 => \N__17640\,
            in3 => \N__19651\,
            lcout => \processor_zipi8.program_counter_i.half_pc_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_0_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17552\,
            lcout => \processor_zipi8.arith_logical_result_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_2_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17530\,
            in1 => \N__18927\,
            in2 => \_gnd_net_\,
            in3 => \N__24167\,
            lcout => OPEN,
            ltout => \processor_zipi8.decode4_strobes_enables_i.un9_flag_enable_type_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_0_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__17519\,
            in1 => \N__23987\,
            in2 => \N__17513\,
            in3 => \N__19943\,
            lcout => OPEN,
            ltout => \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.flag_enable_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__21436\,
            in1 => \N__18928\,
            in2 => \N__17510\,
            in3 => \N__19061\,
            lcout => \processor_zipi8.flag_enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.spm_enable_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__24168\,
            in1 => \N__17483\,
            in2 => \_gnd_net_\,
            in3 => \N__24315\,
            lcout => \processor_zipi8.spm_enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.alu_mux_sel_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000100000"
        )
    port map (
            in0 => \N__19870\,
            in1 => \N__24101\,
            in2 => \N__24341\,
            in3 => \N__21189\,
            lcout => \processor_zipi8.alu_mux_sel_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.use_zero_flag_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__24100\,
            in1 => \N__24333\,
            in2 => \N__21213\,
            in3 => \N__19871\,
            lcout => \processor_zipi8.flags_i.use_zero_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_0_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__33823\,
            in1 => \N__35745\,
            in2 => \N__32230\,
            in3 => \N__31841\,
            lcout => OPEN,
            ltout => \processor_zipi8.alu_result_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNO_3_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18056\,
            in2 => \N__18050\,
            in3 => \N__18043\,
            lcout => \processor_zipi8.flags_i.zero_flag_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNITLO51_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001011010"
        )
    port map (
            in0 => \N__18042\,
            in1 => \N__17974\,
            in2 => \N__19917\,
            in3 => \N__24099\,
            lcout => \processor_zipi8.N_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_1_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__33824\,
            in1 => \N__39127\,
            in2 => \N__39575\,
            in3 => \N__35746\,
            lcout => \processor_zipi8.alu_result_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.arith_logical_sel_1_0_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110110101011"
        )
    port map (
            in0 => \N__24098\,
            in1 => \N__24332\,
            in2 => \N__21212\,
            in3 => \N__19869\,
            lcout => \processor_zipi8.arith_logical_sel_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_2_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__33869\,
            in1 => \N__38310\,
            in2 => \N__38879\,
            in3 => \N__36102\,
            lcout => OPEN,
            ltout => \processor_zipi8.alu_result_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.zero_flag_RNO_2_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20111\,
            in1 => \N__17918\,
            in2 => \N__17912\,
            in3 => \N__17909\,
            lcout => \processor_zipi8.flags_i.zero_flag_3_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__7_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34568\,
            in1 => \N__36668\,
            in2 => \N__33341\,
            in3 => \N__33015\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33680\,
            ce => \N__23437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__7_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34567\,
            in1 => \N__32980\,
            in2 => \N__36627\,
            in3 => \N__33310\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33669\,
            ce => \N__22930\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__7_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34570\,
            in1 => \N__32979\,
            in2 => \N__36803\,
            in3 => \N__33358\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33663\,
            ce => \N__22339\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe12_0_a2_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20848\,
            in1 => \N__22255\,
            in2 => \N__23107\,
            in3 => \N__27392\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe20_0_a2_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27390\,
            in1 => \N__23099\,
            in2 => \N__22290\,
            in3 => \N__20850\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20852\,
            in1 => \N__22266\,
            in2 => \N__23108\,
            in3 => \N__27394\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe4_0_a2_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27389\,
            in1 => \N__23103\,
            in2 => \N__22288\,
            in3 => \N__20847\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20846\,
            in1 => \N__22251\,
            in2 => \N__23165\,
            in3 => \N__27388\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe21_0_a2_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27391\,
            in1 => \N__20534\,
            in2 => \N__22289\,
            in3 => \N__20849\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe6_0_a2_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__23104\,
            in1 => \N__22262\,
            in2 => \N__27460\,
            in3 => \N__20645\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe5_0_a2_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27393\,
            in1 => \N__20535\,
            in2 => \N__22291\,
            in3 => \N__20851\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNINMK21_3_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30835\,
            in1 => \N__18208\,
            in2 => \N__31743\,
            in3 => \N__18194\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_bm_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI1QV11_3_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__18161\,
            in1 => \N__18173\,
            in2 => \N__31693\,
            in3 => \N__30834\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_am_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_3_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18484\,
            in1 => \N__18520\,
            in2 => \_gnd_net_\,
            in3 => \N__37083\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_3_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__18146\,
            in1 => \N__28599\,
            in2 => \N__18212\,
            in3 => \N__28924\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_3_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18209\,
            in1 => \N__18193\,
            in2 => \_gnd_net_\,
            in3 => \N__37084\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_3_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__18089\,
            in1 => \N__18182\,
            in2 => \N__18176\,
            in3 => \N__28600\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_3_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18172\,
            in1 => \N__18160\,
            in2 => \_gnd_net_\,
            in3 => \N__37082\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIHGK21_0_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__18140\,
            in1 => \N__31718\,
            in2 => \N__18122\,
            in3 => \N__30833\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_5_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37299\,
            in1 => \N__18307\,
            in2 => \_gnd_net_\,
            in3 => \N__18325\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_3_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18349\,
            in1 => \N__18340\,
            in2 => \_gnd_net_\,
            in3 => \N__37298\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNILKK21_2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__30973\,
            in1 => \N__18371\,
            in2 => \N__18386\,
            in3 => \N__31581\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI0ESR1_2_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31582\,
            in1 => \N__18461\,
            in2 => \N__18389\,
            in3 => \N__18446\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI0ESR1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_2_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37297\,
            in1 => \N__18382\,
            in2 => \_gnd_net_\,
            in3 => \N__18370\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI4ISR1_3_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100100110001"
        )
    port map (
            in0 => \N__31583\,
            in1 => \N__18359\,
            in2 => \N__18353\,
            in3 => \N__18341\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI4ISR1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIRQK21_5_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__30974\,
            in1 => \N__31584\,
            in2 => \N__18329\,
            in3 => \N__18308\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNICQSR1_5_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31585\,
            in1 => \N__18295\,
            in2 => \N__18281\,
            in3 => \N__18278\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_2_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18226\,
            in1 => \N__18244\,
            in2 => \_gnd_net_\,
            in3 => \N__37294\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIVNV11_2_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__18245\,
            in1 => \N__31390\,
            in2 => \N__18230\,
            in3 => \N__30975\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI2HMP1_2_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__31391\,
            in1 => \N__18557\,
            in2 => \N__18215\,
            in3 => \N__18571\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI2HMP1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_2_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37296\,
            in1 => \_gnd_net_\,
            in2 => \N__18572\,
            in3 => \N__18556\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_2_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__18539\,
            in1 => \N__28544\,
            in2 => \N__18533\,
            in3 => \N__28955\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_2_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28545\,
            in1 => \N__18425\,
            in2 => \N__18530\,
            in3 => \N__18527\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI6LMP1_3_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31392\,
            in1 => \N__18521\,
            in2 => \N__18497\,
            in3 => \N__18485\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI6LMP1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_2_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37295\,
            in1 => \N__18457\,
            in2 => \_gnd_net_\,
            in3 => \N__18445\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIPOK21_4_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__31575\,
            in1 => \N__18409\,
            in2 => \N__30942\,
            in3 => \N__18419\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_4_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__18418\,
            in1 => \N__28957\,
            in2 => \N__18410\,
            in3 => \N__37327\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_4_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28958\,
            in1 => \N__18634\,
            in2 => \N__18392\,
            in3 => \N__18611\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_4_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__18700\,
            in1 => \N__18734\,
            in2 => \N__18686\,
            in3 => \N__28959\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_4_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18743\,
            in2 => \N__18737\,
            in3 => \N__28598\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_4_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__18715\,
            in1 => \N__28956\,
            in2 => \N__37385\,
            in3 => \N__18724\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI3SV11_4_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__31576\,
            in1 => \N__31004\,
            in2 => \N__18728\,
            in3 => \N__18716\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIAPMP1_4_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__18701\,
            in1 => \N__18685\,
            in2 => \N__18665\,
            in3 => \N__31577\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIAPMP1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_4_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35983\,
            in1 => \N__18662\,
            in2 => \_gnd_net_\,
            in3 => \N__18650\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267\,
            ltout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__4_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__35340\,
            in1 => \N__34495\,
            in2 => \N__18638\,
            in3 => \N__35984\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33639\,
            ce => \N__20287\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI8MSR1_4_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31712\,
            in1 => \N__18635\,
            in2 => \N__18620\,
            in3 => \N__18610\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI8MSR1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_1_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18596\,
            in1 => \N__18584\,
            in2 => \_gnd_net_\,
            in3 => \N__35982\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198\,
            ltout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34494\,
            in1 => \N__36850\,
            in2 => \N__19106\,
            in3 => \N__39494\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33639\,
            ce => \N__20287\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIS9SR1_1_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__20753\,
            in1 => \N__20732\,
            in2 => \N__20951\,
            in3 => \N__31708\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI1P541_4_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30917\,
            in1 => \N__24953\,
            in2 => \N__31741\,
            in3 => \N__25109\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_4_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24952\,
            in1 => \N__25108\,
            in2 => \_gnd_net_\,
            in3 => \N__37429\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_3_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19103\,
            in2 => \_gnd_net_\,
            in3 => \N__19085\,
            lcout => \processor_zipi8.arith_logical_result_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001010"
        )
    port map (
            in0 => \N__18925\,
            in1 => \N__19963\,
            in2 => \N__19079\,
            in3 => \N__24166\,
            lcout => OPEN,
            ltout => \processor_zipi8.decode4_strobes_enables_i.register_enable_type_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.register_enable_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__21391\,
            in1 => \N__19031\,
            in2 => \N__18935\,
            in3 => \N__18926\,
            lcout => \processor_zipi8.register_enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__18812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19258\,
            lcout => \processor_zipi8.arith_logical_result_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical4_process_carry_arith_logical_28_4_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__19776\,
            in1 => \N__21846\,
            in2 => \N__19259\,
            in3 => \N__18811\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4\,
            ltout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical5_process_carry_arith_logical_34_5_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__18797\,
            in1 => \N__19321\,
            in2 => \N__19334\,
            in3 => \N__19777\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_34_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_5_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__19322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19310\,
            lcout => \processor_zipi8.arith_logical_result_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.flags_i.carry_flag_RNO_6_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35297\,
            in1 => \N__37899\,
            in2 => \N__38731\,
            in3 => \N__30207\,
            lcout => \processor_zipi8.flags_i.parity_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000101"
        )
    port map (
            in0 => \N__21683\,
            in1 => \N__23989\,
            in2 => \N__19556\,
            in3 => \N__19499\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__19397\,
            in1 => \N__21684\,
            in2 => \N__19298\,
            in3 => \N__19295\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tz_4_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110111111"
        )
    port map (
            in0 => \N__19203\,
            in1 => \N__21821\,
            in2 => \N__19782\,
            in3 => \N__19472\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tzZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_4_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000000010"
        )
    port map (
            in0 => \N__23990\,
            in1 => \N__19234\,
            in2 => \N__21836\,
            in3 => \N__19536\,
            lcout => OPEN,
            ltout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__19236\,
            in1 => \N__19268\,
            in2 => \N__19262\,
            in3 => \N__19112\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_4_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001101111111"
        )
    port map (
            in0 => \N__19471\,
            in1 => \N__19235\,
            in2 => \N__21835\,
            in3 => \N__19204\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001011111"
        )
    port map (
            in0 => \N__21682\,
            in1 => \N__19617\,
            in2 => \N__19555\,
            in3 => \N__21546\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_1_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110111011101"
        )
    port map (
            in0 => \N__21547\,
            in1 => \N__19493\,
            in2 => \N__19482\,
            in3 => \N__19751\,
            lcout => \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNINIG61_4_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__31009\,
            in1 => \N__19376\,
            in2 => \N__32528\,
            in3 => \N__31573\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI4AK32_4_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31574\,
            in1 => \N__23359\,
            in2 => \N__19391\,
            in3 => \N__33731\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI4AK32_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_4_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37424\,
            in1 => \N__22978\,
            in2 => \_gnd_net_\,
            in3 => \N__27707\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_4_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__28647\,
            in1 => \N__19388\,
            in2 => \N__19379\,
            in3 => \N__29001\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_4_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37425\,
            in1 => \_gnd_net_\,
            in2 => \N__23360\,
            in3 => \N__33730\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_4_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19375\,
            in1 => \N__32524\,
            in2 => \_gnd_net_\,
            in3 => \N__37426\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_4_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__19358\,
            in1 => \N__19352\,
            in2 => \N__19346\,
            in3 => \N__28648\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_4_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__25603\,
            in1 => \N__19979\,
            in2 => \N__25160\,
            in3 => \N__25763\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4alu_i.arith_logical_sel_1_2_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__19918\,
            in1 => \N__24310\,
            in2 => \_gnd_net_\,
            in3 => \N__24126\,
            lcout => \processor_zipi8.arith_logical_sel_1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_3_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__28646\,
            in1 => \N__23579\,
            in2 => \N__20153\,
            in3 => \N__19664\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_3_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__25601\,
            in1 => \N__19682\,
            in2 => \N__19670\,
            in3 => \N__25762\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_3_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21931\,
            in1 => \N__23485\,
            in2 => \_gnd_net_\,
            in3 => \N__37423\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_3_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__25970\,
            in1 => \N__28645\,
            in2 => \N__19667\,
            in3 => \N__28997\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_3_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__27821\,
            in1 => \N__25602\,
            in2 => \N__26267\,
            in3 => \N__19658\,
            lcout => \processor_zipi8.sy_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIPPE01_3_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__31008\,
            in1 => \N__23600\,
            in2 => \N__23621\,
            in3 => \N__31572\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_bm_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI8OGN1_3_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__20165\,
            in1 => \N__22388\,
            in2 => \N__19643\,
            in3 => \N__31570\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI8OGN1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU6AG4_3_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__20099\,
            in1 => \N__27312\,
            in2 => \N__20105\,
            in3 => \N__27609\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIHPTE1_3_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__21932\,
            in1 => \N__31569\,
            in2 => \N__23486\,
            in3 => \N__31007\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_am_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIONE42_3_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26207\,
            in1 => \N__25985\,
            in2 => \N__20102\,
            in3 => \N__31571\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIONE42_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINP2G8_3_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__27313\,
            in1 => \N__20093\,
            in2 => \N__20081\,
            in3 => \N__20066\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINP2G8_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5OSHH_3_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__22169\,
            in1 => \N__27110\,
            in2 => \N__20060\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.sx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__0_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35976\,
            in1 => \N__33903\,
            in2 => \N__32289\,
            in3 => \N__31997\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33679\,
            ce => \N__20140\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__1_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__33902\,
            in1 => \N__39544\,
            in2 => \N__39227\,
            in3 => \N__35981\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33679\,
            ce => \N__20140\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__2_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__35977\,
            in1 => \N__38847\,
            in2 => \N__34276\,
            in3 => \N__38446\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33679\,
            ce => \N__20140\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_2_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22399\,
            in1 => \N__21790\,
            in2 => \_gnd_net_\,
            in3 => \N__37503\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__3_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35978\,
            in1 => \N__33904\,
            in2 => \N__38159\,
            in3 => \N__37627\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33679\,
            ce => \N__20140\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_3_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22387\,
            in1 => \N__20164\,
            in2 => \_gnd_net_\,
            in3 => \N__37504\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__4_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__35979\,
            in1 => \N__35347\,
            in2 => \N__35097\,
            in3 => \N__33908\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33679\,
            ce => \N__20140\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__5_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__30089\,
            in1 => \N__35980\,
            in2 => \N__34078\,
            in3 => \N__30390\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33679\,
            ce => \N__20140\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_4_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__33825\,
            in1 => \N__35007\,
            in2 => \N__35413\,
            in3 => \N__36101\,
            lcout => \processor_zipi8.alu_result_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__7_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34325\,
            in1 => \N__33002\,
            in2 => \N__36792\,
            in3 => \N__33327\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33690\,
            ce => \N__27781\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__5_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__30464\,
            in1 => \N__34580\,
            in2 => \N__30134\,
            in3 => \N__36625\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33682\,
            ce => \N__32497\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__6_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34579\,
            in1 => \N__36623\,
            in2 => \N__29782\,
            in3 => \N__29291\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33682\,
            ce => \N__32497\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__7_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__33301\,
            in1 => \N__36624\,
            in2 => \N__33010\,
            in3 => \N__34581\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33682\,
            ce => \N__32497\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI7V541_7_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__20186\,
            in1 => \N__31734\,
            in2 => \N__31022\,
            in3 => \N__21581\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI43VU1_7_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31735\,
            in1 => \N__20203\,
            in2 => \N__20237\,
            in3 => \N__22577\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI43VU1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNITOG61_7_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__21607\,
            in1 => \N__31736\,
            in2 => \N__32714\,
            in3 => \N__31013\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIGMK32_7_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31737\,
            in1 => \N__23315\,
            in2 => \N__20234\,
            in3 => \N__23872\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIGMK32_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIGUM4_7_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__20231\,
            in1 => \N__27286\,
            in2 => \N__20225\,
            in3 => \N__27629\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_7_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20204\,
            in1 => \N__22576\,
            in2 => \_gnd_net_\,
            in3 => \N__37355\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_7_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__20171\,
            in1 => \N__28658\,
            in2 => \N__20189\,
            in3 => \N__28968\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_7_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21580\,
            in1 => \N__20185\,
            in2 => \_gnd_net_\,
            in3 => \N__37354\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe31_0_a2_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20642\,
            in1 => \N__22268\,
            in2 => \N__20541\,
            in3 => \N__27430\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe19_0_a2_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27428\,
            in1 => \N__20332\,
            in2 => \N__22292\,
            in3 => \N__20639\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe7_0_a2_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20644\,
            in1 => \N__22267\,
            in2 => \N__20542\,
            in3 => \N__27429\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe3_0_a2_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27433\,
            in1 => \N__20333\,
            in2 => \N__22294\,
            in3 => \N__20643\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe14_0_a2_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20638\,
            in1 => \N__22279\,
            in2 => \N__23105\,
            in3 => \N__27435\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe22_0_a2_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27432\,
            in1 => \N__23092\,
            in2 => \N__22293\,
            in3 => \N__20640\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe30_0_a2_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20641\,
            in1 => \N__22272\,
            in2 => \N__23106\,
            in3 => \N__27431\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27434\,
            in1 => \N__20527\,
            in2 => \N__22295\,
            in3 => \N__20853\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI7JI91_4_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30822\,
            in1 => \N__26075\,
            in2 => \N__31703\,
            in3 => \N__24521\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNII4IQ1_4_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__24482\,
            in1 => \N__24499\,
            in2 => \N__20258\,
            in3 => \N__31623\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNII4IQ1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNI12F01_7_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30823\,
            in1 => \N__20489\,
            in2 => \N__31704\,
            in3 => \N__20468\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIO8HN1_7_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__20440\,
            in1 => \N__20426\,
            in2 => \N__20255\,
            in3 => \N__31624\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIO8HN1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_7_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20485\,
            in1 => \N__20467\,
            in2 => \_gnd_net_\,
            in3 => \N__37214\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_7_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37215\,
            in1 => \_gnd_net_\,
            in2 => \N__20441\,
            in3 => \N__20425\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIJJE01_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__31616\,
            in1 => \N__23276\,
            in2 => \N__30921\,
            in3 => \N__23411\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe24_0_a2_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20831\,
            in1 => \N__27289\,
            in2 => \N__22283\,
            in3 => \N__23146\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_5_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37332\,
            in1 => \N__29812\,
            in2 => \_gnd_net_\,
            in3 => \N__22648\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_5_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__20339\,
            in1 => \N__20666\,
            in2 => \N__20402\,
            in3 => \N__28602\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIO5SR1_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__20386\,
            in1 => \N__20369\,
            in2 => \N__20348\,
            in3 => \N__31713\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIO5SR1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_5_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22948\,
            in1 => \N__22747\,
            in2 => \_gnd_net_\,
            in3 => \N__37328\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_5_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37330\,
            in1 => \N__23338\,
            in2 => \_gnd_net_\,
            in3 => \N__23890\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_5_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22768\,
            in1 => \N__24940\,
            in2 => \_gnd_net_\,
            in3 => \N__37329\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_5_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__28601\,
            in1 => \N__20675\,
            in2 => \N__20669\,
            in3 => \N__28885\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_6_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29095\,
            in1 => \N__22442\,
            in2 => \_gnd_net_\,
            in3 => \N__37331\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_2_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20873\,
            in2 => \_gnd_net_\,
            in3 => \N__31428\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIBJTE1_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__31425\,
            in1 => \N__23534\,
            in2 => \N__31017\,
            in3 => \N__21979\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNICBE42_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__25448\,
            in1 => \N__25913\,
            in2 => \N__20582\,
            in3 => \N__31426\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNICBE42_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6E9G4_0_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__27287\,
            in1 => \N__27594\,
            in2 => \N__20579\,
            in3 => \N__20768\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI781G8_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__27288\,
            in1 => \N__20576\,
            in2 => \N__20564\,
            in3 => \N__20561\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI781G8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27595\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20872\,
            in2 => \_gnd_net_\,
            in3 => \N__31427\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNISBGN1_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__31424\,
            in1 => \N__20900\,
            in2 => \N__21920\,
            in3 => \N__20777\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNISBGN1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIUCMP1_1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31707\,
            in1 => \N__21017\,
            in2 => \N__20762\,
            in3 => \N__20999\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNITLV11_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__20714\,
            in1 => \N__31706\,
            in2 => \N__20696\,
            in3 => \N__30848\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__37323\,
            in1 => \N__20965\,
            in2 => \N__28998\,
            in3 => \N__20980\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__20752\,
            in1 => \N__20731\,
            in2 => \N__20720\,
            in3 => \N__28954\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20987\,
            in2 => \N__20717\,
            in3 => \N__28587\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_1_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__20713\,
            in1 => \N__28949\,
            in2 => \N__20695\,
            in3 => \N__37322\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28950\,
            in1 => \N__21016\,
            in2 => \N__21002\,
            in3 => \N__20998\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIJIK21_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__20981\,
            in1 => \N__31705\,
            in2 => \N__20969\,
            in3 => \N__30847\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_7_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010101"
        )
    port map (
            in0 => \N__20942\,
            in1 => \N__21587\,
            in2 => \N__20912\,
            in3 => \N__28586\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__28927\,
            in1 => \N__37301\,
            in2 => \N__21980\,
            in3 => \N__23533\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28929\,
            in1 => \N__25912\,
            in2 => \N__20918\,
            in3 => \N__25447\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_0_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__28585\,
            in1 => \_gnd_net_\,
            in2 => \N__20915\,
            in3 => \N__20879\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_7_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37303\,
            in1 => \N__23311\,
            in2 => \_gnd_net_\,
            in3 => \N__23873\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_0_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__28926\,
            in1 => \N__37300\,
            in2 => \N__23275\,
            in3 => \N__23407\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_0_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28928\,
            in1 => \N__21913\,
            in2 => \N__20903\,
            in3 => \N__20896\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_7_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32701\,
            in1 => \N__21608\,
            in2 => \_gnd_net_\,
            in3 => \N__37302\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__5_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__30034\,
            in1 => \N__36525\,
            in2 => \N__34824\,
            in3 => \N__30269\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33650\,
            ce => \N__25091\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__6_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36524\,
            in1 => \N__29642\,
            in2 => \N__29397\,
            in3 => \N__34711\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33650\,
            ce => \N__25091\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__7_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__32823\,
            in1 => \N__36526\,
            in2 => \N__34825\,
            in3 => \N__33219\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33650\,
            ce => \N__25091\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_6_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21507\,
            in1 => \N__21389\,
            in2 => \_gnd_net_\,
            in3 => \N__23191\,
            lcout => \processor_zipi8.port_id_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI7UF21_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21388\,
            in1 => \N__21533\,
            in2 => \_gnd_net_\,
            in3 => \N__21508\,
            lcout => \processor_zipi8.pc_vector_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIC1G21_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21470\,
            in1 => \N__21390\,
            in2 => \_gnd_net_\,
            in3 => \N__37427\,
            lcout => \processor_zipi8.pc_vector_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.sel_of_out_port_value_i.un1_sx_7_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37428\,
            in1 => \N__21226\,
            in2 => \_gnd_net_\,
            in3 => \N__21110\,
            lcout => \LED1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNILLE01_1_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30945\,
            in1 => \N__25405\,
            in2 => \N__31568\,
            in3 => \N__25424\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI0GGN1_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__25370\,
            in1 => \N__25391\,
            in2 => \N__21755\,
            in3 => \N__31398\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_119_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIEM9G4_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__27277\,
            in1 => \N__21746\,
            in2 => \N__21752\,
            in3 => \N__27564\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIDLTE1_1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23249\,
            in1 => \N__31393\,
            in2 => \N__23510\,
            in3 => \N__30944\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIGFE42_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31394\,
            in1 => \N__25883\,
            in2 => \N__21749\,
            in3 => \N__26033\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINO1G8_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__21740\,
            in1 => \N__27278\,
            in2 => \N__21731\,
            in3 => \N__21716\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5MQHH_1_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__22159\,
            in1 => \_gnd_net_\,
            in2 => \N__21710\,
            in3 => \N__26477\,
            lcout => \processor_zipi8.sx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFIBI8_4_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__26666\,
            in1 => \N__21614\,
            in2 => \N__21650\,
            in3 => \N__27275\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFIBI8_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIOMUU1_4_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__22979\,
            in1 => \N__27706\,
            in2 => \N__21638\,
            in3 => \N__31688\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIOMUU1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQNTM4_4_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__21623\,
            in1 => \N__27273\,
            in2 => \N__21617\,
            in3 => \N__27610\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7A3G8_4_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__27276\,
            in1 => \N__21896\,
            in2 => \N__21884\,
            in3 => \N__21803\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7A3G8_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5PTHH_4_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21869\,
            in2 => \N__21863\,
            in3 => \N__22231\,
            lcout => \processor_zipi8.sx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNISRE42_4_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26189\,
            in1 => \N__25283\,
            in2 => \N__25121\,
            in3 => \N__31689\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNISRE42_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6FAG4_4_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__23177\,
            in1 => \N__27274\,
            in2 => \N__21806\,
            in3 => \N__27611\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIFNTE1_2_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25489\,
            in1 => \N__31512\,
            in2 => \N__25508\,
            in3 => \N__31006\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNINNE01_2_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__31005\,
            in1 => \N__23387\,
            in2 => \N__31673\,
            in3 => \N__23375\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI4KGN1_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__22403\,
            in1 => \N__21797\,
            in2 => \N__21779\,
            in3 => \N__31513\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI4KGN1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIKJE42_2_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31514\,
            in1 => \N__25859\,
            in2 => \N__21776\,
            in3 => \N__26009\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIKJE42_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMU9G4_2_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__21767\,
            in1 => \N__27314\,
            in2 => \N__21758\,
            in3 => \N__27605\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI792G8_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__27315\,
            in1 => \N__22328\,
            in2 => \N__22313\,
            in3 => \N__22310\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI792G8_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5NRHH_2_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__22230\,
            in1 => \_gnd_net_\,
            in2 => \N__22052\,
            in3 => \N__27041\,
            lcout => \processor_zipi8.sx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__0_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34826\,
            in1 => \N__32264\,
            in2 => \N__32027\,
            in3 => \N__35847\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33681\,
            ce => \N__25346\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__2_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__35844\,
            in1 => \N__38830\,
            in2 => \N__38506\,
            in3 => \N__34828\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33681\,
            ce => \N__25346\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_3_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21962\,
            in1 => \N__21950\,
            in2 => \_gnd_net_\,
            in3 => \N__35843\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266\,
            ltout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__3_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__35845\,
            in1 => \N__38071\,
            in2 => \N__21935\,
            in3 => \N__34830\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33681\,
            ce => \N__25346\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34827\,
            in1 => \N__39178\,
            in2 => \N__39635\,
            in3 => \N__35848\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33681\,
            ce => \N__25346\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__5_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35846\,
            in1 => \N__34829\,
            in2 => \N__30490\,
            in3 => \N__30024\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33681\,
            ce => \N__25346\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34068\,
            in1 => \N__35973\,
            in2 => \N__32403\,
            in3 => \N__32022\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33689\,
            ce => \N__22352\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35969\,
            in1 => \N__34071\,
            in2 => \N__39644\,
            in3 => \N__39225\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33689\,
            ce => \N__22352\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__2_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34069\,
            in1 => \N__35975\,
            in2 => \N__38518\,
            in3 => \N__38874\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33689\,
            ce => \N__22352\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__3_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__35970\,
            in1 => \N__38144\,
            in2 => \N__37706\,
            in3 => \N__34073\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33689\,
            ce => \N__22352\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__4_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34070\,
            in1 => \N__35974\,
            in2 => \N__35230\,
            in3 => \N__35530\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33689\,
            ce => \N__22352\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__5_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__35971\,
            in1 => \N__30485\,
            in2 => \N__30088\,
            in3 => \N__34074\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33689\,
            ce => \N__22352\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_5_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23704\,
            in1 => \N__23686\,
            in2 => \_gnd_net_\,
            in3 => \N__37487\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__6_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35972\,
            in1 => \N__34072\,
            in2 => \N__29773\,
            in3 => \N__29396\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33689\,
            ce => \N__22352\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__6_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34326\,
            in1 => \N__29447\,
            in2 => \N__36793\,
            in3 => \N__29735\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33701\,
            ce => \N__24413\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__5_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34796\,
            in1 => \N__36656\,
            in2 => \N__30146\,
            in3 => \N__30500\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33692\,
            ce => \N__27679\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__6_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36655\,
            in1 => \N__34798\,
            in2 => \N__29783\,
            in3 => \N__29445\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33692\,
            ce => \N__27679\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__7_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34797\,
            in1 => \N__36657\,
            in2 => \N__33021\,
            in3 => \N__33302\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33692\,
            ce => \N__27679\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_6_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22592\,
            in1 => \N__22609\,
            in2 => \_gnd_net_\,
            in3 => \N__37293\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIRMG61_6_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22438\,
            in1 => \N__31679\,
            in2 => \N__29102\,
            in3 => \N__30981\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNICIK32_6_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31681\,
            in1 => \N__24572\,
            in2 => \N__22424\,
            in3 => \N__24548\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNICIK32_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA8UM4_6_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22625\,
            in1 => \N__27384\,
            in2 => \N__22421\,
            in3 => \N__27628\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFJCI8_6_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__27385\,
            in1 => \N__24362\,
            in2 => \N__22418\,
            in3 => \N__22598\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFJCI8_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI5T541_6_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__24866\,
            in1 => \N__31677\,
            in2 => \N__24890\,
            in3 => \N__30980\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI0VUU1_6_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31678\,
            in1 => \N__22913\,
            in2 => \N__22628\,
            in3 => \N__22897\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI0VUU1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIQCIQ1_6_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110010001"
        )
    port map (
            in0 => \N__23846\,
            in1 => \N__31680\,
            in2 => \N__22619\,
            in3 => \N__22591\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIQCIQ1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__0_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34799\,
            in1 => \N__36666\,
            in2 => \N__32350\,
            in3 => \N__32092\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33671\,
            ce => \N__27774\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__1_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36662\,
            in1 => \N__39596\,
            in2 => \N__39282\,
            in3 => \N__34803\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33671\,
            ce => \N__27774\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__3_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36663\,
            in1 => \N__34801\,
            in2 => \N__38188\,
            in3 => \N__37793\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33671\,
            ce => \N__27774\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__4_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34800\,
            in1 => \N__36667\,
            in2 => \N__35229\,
            in3 => \N__35546\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33671\,
            ce => \N__27774\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__5_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36664\,
            in1 => \N__34802\,
            in2 => \N__30471\,
            in3 => \N__30145\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33671\,
            ce => \N__27774\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_5_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22663\,
            in1 => \N__24424\,
            in2 => \_gnd_net_\,
            in3 => \N__37254\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__6_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36665\,
            in1 => \N__29743\,
            in2 => \N__29370\,
            in3 => \N__34804\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33671\,
            ce => \N__27774\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI1L181_5_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__28037\,
            in1 => \N__30837\,
            in2 => \N__31733\,
            in3 => \N__28216\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_5_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37213\,
            in1 => \_gnd_net_\,
            in2 => \N__28217\,
            in3 => \N__28036\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_5_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__22682\,
            in1 => \N__28575\,
            in2 => \N__22709\,
            in3 => \N__28925\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_5_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28576\,
            in1 => \N__22706\,
            in2 => \N__22700\,
            in3 => \N__22676\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_5_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26443\,
            in1 => \N__29071\,
            in2 => \_gnd_net_\,
            in3 => \N__37211\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_5_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37212\,
            in1 => \_gnd_net_\,
            in2 => \N__24353\,
            in3 => \N__26050\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI9LI91_5_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__26051\,
            in1 => \N__24352\,
            in2 => \N__31732\,
            in3 => \N__30836\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIM8IQ1_5_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__24425\,
            in1 => \N__31663\,
            in2 => \N__22670\,
            in3 => \N__22667\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIPKG61_5_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22652\,
            in1 => \N__31539\,
            in2 => \N__29816\,
            in3 => \N__30910\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI8EK32_5_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31541\,
            in1 => \N__23339\,
            in2 => \N__22631\,
            in3 => \N__23894\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_243_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI20UM4_5_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22730\,
            in1 => \N__27320\,
            in2 => \N__22808\,
            in3 => \N__27632\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV2CI8_5_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__27321\,
            in1 => \N__22805\,
            in2 => \N__22793\,
            in3 => \N__22715\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI3R541_5_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22772\,
            in1 => \N__31537\,
            in2 => \N__24941\,
            in3 => \N__30909\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNISQUU1_5_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31538\,
            in1 => \N__22949\,
            in2 => \N__22751\,
            in3 => \N__22748\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIOEMM1_5_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26444\,
            in1 => \N__29075\,
            in2 => \N__22724\,
            in3 => \N__31540\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34633\,
            in1 => \N__32398\,
            in2 => \N__32100\,
            in3 => \N__36403\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33651\,
            ce => \N__22937\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__39595\,
            in1 => \N__34637\,
            in2 => \N__39290\,
            in3 => \N__36377\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33651\,
            ce => \N__22937\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34634\,
            in1 => \N__36404\,
            in2 => \N__38568\,
            in3 => \N__38799\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33651\,
            ce => \N__22937\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__3_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111000000010"
        )
    port map (
            in0 => \N__38118\,
            in1 => \N__34638\,
            in2 => \N__36605\,
            in3 => \N__37703\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33651\,
            ce => \N__22937\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34635\,
            in1 => \N__36405\,
            in2 => \N__35234\,
            in3 => \N__35472\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33651\,
            ce => \N__22937\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__5_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__30069\,
            in1 => \N__34639\,
            in2 => \N__36606\,
            in3 => \N__30489\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33651\,
            ce => \N__22937\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__6_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34636\,
            in1 => \N__36406\,
            in2 => \N__29406\,
            in3 => \N__29722\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33651\,
            ce => \N__22937\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_6_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22909\,
            in1 => \N__22898\,
            in2 => \_gnd_net_\,
            in3 => \N__37356\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIUGIQ1_7_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__22817\,
            in1 => \N__30566\,
            in2 => \N__22838\,
            in3 => \N__31684\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIUGIQ1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_7_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22868\,
            in1 => \N__22856\,
            in2 => \_gnd_net_\,
            in3 => \N__36143\,
            lcout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269\,
            ltout => \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36144\,
            in1 => \N__33203\,
            in2 => \N__22841\,
            in3 => \N__34467\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33640\,
            ce => \N__24409\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_7_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37372\,
            in1 => \N__22834\,
            in2 => \_gnd_net_\,
            in3 => \N__22816\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIRRE01_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25259\,
            in1 => \N__31682\,
            in2 => \N__25241\,
            in3 => \N__30898\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNICSGN1_4_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31683\,
            in1 => \N__25220\,
            in2 => \N__23180\,
            in3 => \N__25196\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNICSGN1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27590\,
            in2 => \_gnd_net_\,
            in3 => \N__30899\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__30900\,
            in1 => \_gnd_net_\,
            in2 => \N__27624\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__27001\,
            in1 => \N__23255\,
            in2 => \N__24815\,
            in3 => \N__28933\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28556\,
            in2 => \N__23057\,
            in3 => \N__23051\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_1_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__30553\,
            in1 => \N__28931\,
            in2 => \N__32650\,
            in3 => \N__37441\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28932\,
            in1 => \N__24760\,
            in2 => \N__23054\,
            in3 => \N__31801\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__25635\,
            in1 => \N__25737\,
            in2 => \N__23045\,
            in3 => \N__23027\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25636\,
            in1 => \N__24689\,
            in2 => \N__23021\,
            in3 => \N__23018\,
            lcout => \processor_zipi8.sy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_1_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__24719\,
            in1 => \N__28930\,
            in2 => \N__24832\,
            in3 => \N__37440\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25061\,
            in1 => \N__26552\,
            in2 => \_gnd_net_\,
            in3 => \N__28558\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23248\,
            in1 => \N__28999\,
            in2 => \N__23509\,
            in3 => \N__37451\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29000\,
            in1 => \N__25882\,
            in2 => \N__23231\,
            in3 => \N__26032\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__28557\,
            in1 => \_gnd_net_\,
            in2 => \N__23228\,
            in3 => \N__25352\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__25638\,
            in1 => \N__23225\,
            in2 => \N__23216\,
            in3 => \N__25755\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__28559\,
            in1 => \N__32594\,
            in2 => \N__38909\,
            in3 => \N__24959\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__25639\,
            in1 => \N__23213\,
            in2 => \N__23207\,
            in3 => \N__23204\,
            lcout => \processor_zipi8.sy_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34190\,
            in1 => \N__32362\,
            in2 => \N__32109\,
            in3 => \N__36192\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36186\,
            in1 => \N__39450\,
            in2 => \N__39260\,
            in3 => \N__34196\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34191\,
            in1 => \N__36190\,
            in2 => \N__38552\,
            in3 => \N__38878\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36187\,
            in1 => \N__34194\,
            in2 => \N__38145\,
            in3 => \N__37661\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__4_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__36191\,
            in2 => \N__35535\,
            in3 => \N__35123\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__5_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36188\,
            in1 => \N__30439\,
            in2 => \N__30090\,
            in3 => \N__34197\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__6_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34193\,
            in1 => \N__29393\,
            in2 => \N__29780\,
            in3 => \N__36193\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__7_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36189\,
            in1 => \N__34195\,
            in2 => \N__33294\,
            in3 => \N__32792\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33664\,
            ce => \N__23291\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36279\,
            in1 => \N__34183\,
            in2 => \N__32437\,
            in3 => \N__32079\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33670\,
            ce => \N__23438\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__39198\,
            in1 => \N__39535\,
            in2 => \N__34468\,
            in3 => \N__36284\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33670\,
            ce => \N__23438\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36280\,
            in1 => \N__38834\,
            in2 => \N__38530\,
            in3 => \N__34187\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33670\,
            ce => \N__23438\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34180\,
            in1 => \N__36282\,
            in2 => \N__37704\,
            in3 => \N__38078\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33670\,
            ce => \N__23438\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__4_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__36281\,
            in1 => \N__35145\,
            in2 => \N__35556\,
            in3 => \N__34188\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33670\,
            ce => \N__23438\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34181\,
            in1 => \N__30067\,
            in2 => \N__36523\,
            in3 => \N__30440\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33670\,
            ce => \N__23438\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_5_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23722\,
            in1 => \N__23743\,
            in2 => \_gnd_net_\,
            in3 => \N__37505\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__6_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34182\,
            in1 => \N__36283\,
            in2 => \N__29407\,
            in3 => \N__29764\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33670\,
            ce => \N__23438\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34818\,
            in1 => \N__32323\,
            in2 => \N__32080\,
            in3 => \N__36142\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33683\,
            ce => \N__23570\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36137\,
            in1 => \N__39568\,
            in2 => \N__39248\,
            in3 => \N__34823\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33683\,
            ce => \N__23570\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34819\,
            in1 => \N__36139\,
            in2 => \N__38461\,
            in3 => \N__38835\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33683\,
            ce => \N__23570\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23386\,
            in1 => \N__23371\,
            in2 => \_gnd_net_\,
            in3 => \N__37488\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__3_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34820\,
            in1 => \N__36140\,
            in2 => \N__37668\,
            in3 => \N__38079\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33683\,
            ce => \N__23570\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__23611\,
            in1 => \_gnd_net_\,
            in2 => \N__23596\,
            in3 => \N__37489\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__4_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34821\,
            in1 => \N__36141\,
            in2 => \N__35204\,
            in3 => \N__35521\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33683\,
            ce => \N__23570\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__5_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36138\,
            in1 => \N__34822\,
            in2 => \N__30491\,
            in3 => \N__30115\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33683\,
            ce => \N__23570\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34810\,
            in1 => \N__35880\,
            in2 => \N__32316\,
            in3 => \N__31958\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35876\,
            in1 => \N__34814\,
            in2 => \N__39643\,
            in3 => \N__39240\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34811\,
            in1 => \N__35881\,
            in2 => \N__38517\,
            in3 => \N__38836\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35877\,
            in1 => \N__34815\,
            in2 => \N__38146\,
            in3 => \N__37654\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34812\,
            in1 => \N__35882\,
            in2 => \N__35231\,
            in3 => \N__35523\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__5_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35878\,
            in1 => \N__34816\,
            in2 => \N__30509\,
            in3 => \N__30116\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__6_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34813\,
            in1 => \N__35883\,
            in2 => \N__29408\,
            in3 => \N__29781\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__7_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35879\,
            in1 => \N__34817\,
            in2 => \N__33335\,
            in3 => \N__32793\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33691\,
            ce => \N__23762\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNITTE01_5_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23747\,
            in1 => \N__31612\,
            in2 => \N__23732\,
            in3 => \N__30982\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIG0HN1_5_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31613\,
            in1 => \N__23711\,
            in2 => \N__23693\,
            in3 => \N__23690\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNILTTE1_5_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25048\,
            in1 => \N__31614\,
            in2 => \N__25033\,
            in3 => \N__30983\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI00F42_5_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31615\,
            in1 => \N__26126\,
            in2 => \N__23675\,
            in3 => \N__26114\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIENAG4_5_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__23672\,
            in1 => \N__27285\,
            in2 => \N__23666\,
            in3 => \N__27630\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.x12_bit_program_address_generator_i.return_vector_3_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23648\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.decode4_strobes_enables_i.un29_flag_enable_type_0_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24337\,
            in2 => \_gnd_net_\,
            in3 => \N__24111\,
            lcout => \processor_zipi8.un28_carry_flag_value_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__4_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36315\,
            in1 => \N__34189\,
            in2 => \N__35567\,
            in3 => \N__35203\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33704\,
            ce => \N__25958\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__5_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34881\,
            in1 => \N__36659\,
            in2 => \N__30155\,
            in3 => \N__30493\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33703\,
            ce => \N__33385\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__6_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36658\,
            in1 => \N__29771\,
            in2 => \N__29446\,
            in3 => \N__34883\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33703\,
            ce => \N__33385\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__7_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34882\,
            in1 => \N__36660\,
            in2 => \N__33011\,
            in3 => \N__33339\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33703\,
            ce => \N__33385\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIBNI91_6_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__31674\,
            in1 => \N__26315\,
            in2 => \N__24449\,
            in3 => \N__30845\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_6_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37136\,
            in1 => \N__28198\,
            in2 => \_gnd_net_\,
            in3 => \N__28018\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_6_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__24377\,
            in1 => \N__28640\,
            in2 => \N__23840\,
            in3 => \N__28973\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_6_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28641\,
            in1 => \N__23837\,
            in2 => \N__23831\,
            in3 => \N__24371\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_6_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26419\,
            in1 => \N__29053\,
            in2 => \_gnd_net_\,
            in3 => \N__37134\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_6_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37135\,
            in1 => \N__26314\,
            in2 => \_gnd_net_\,
            in3 => \N__24445\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI3N181_6_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__31675\,
            in1 => \N__28199\,
            in2 => \N__28022\,
            in3 => \N__30846\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNISIMM1_6_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__29054\,
            in1 => \N__26420\,
            in2 => \N__24365\,
            in3 => \N__31676\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNISIMM1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34842\,
            in1 => \N__36612\,
            in2 => \N__32351\,
            in3 => \N__32093\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__1_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36608\,
            in1 => \N__39630\,
            in2 => \N__39283\,
            in3 => \N__34851\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34843\,
            in1 => \N__36613\,
            in2 => \N__38567\,
            in3 => \N__38820\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36609\,
            in1 => \N__34845\,
            in2 => \N__38189\,
            in3 => \N__37754\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__4_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__35228\,
            in1 => \N__35494\,
            in2 => \N__34880\,
            in3 => \N__36849\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__5_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36610\,
            in1 => \N__34846\,
            in2 => \N__30472\,
            in3 => \N__30144\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__6_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34844\,
            in1 => \N__36614\,
            in2 => \N__29369\,
            in3 => \N__29744\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__7_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36611\,
            in1 => \N__33338\,
            in2 => \N__33028\,
            in3 => \N__34850\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33685\,
            ce => \N__24437\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34618\,
            in1 => \N__36796\,
            in2 => \N__32439\,
            in3 => \N__32121\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33672\,
            ce => \N__24408\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24631\,
            in1 => \N__24652\,
            in2 => \_gnd_net_\,
            in3 => \N__37216\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__1_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34619\,
            in1 => \N__39631\,
            in2 => \N__39229\,
            in3 => \N__36799\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33672\,
            ce => \N__24408\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__2_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__36794\,
            in1 => \N__38533\,
            in2 => \N__38891\,
            in3 => \N__34624\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33672\,
            ce => \N__24408\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__3_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34620\,
            in1 => \N__36797\,
            in2 => \N__38187\,
            in3 => \N__37753\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33672\,
            ce => \N__24408\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_3_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26383\,
            in1 => \N__26365\,
            in2 => \_gnd_net_\,
            in3 => \N__37217\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__4_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__35093\,
            in1 => \N__36798\,
            in2 => \N__34795\,
            in3 => \N__35547\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33672\,
            ce => \N__24408\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36795\,
            in1 => \N__30448\,
            in2 => \N__30121\,
            in3 => \N__34625\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33672\,
            ce => \N__24408\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_6_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010101"
        )
    port map (
            in0 => \N__24455\,
            in1 => \N__24620\,
            in2 => \N__24530\,
            in3 => \N__28442\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_4_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__28060\,
            in1 => \N__28780\,
            in2 => \N__28240\,
            in3 => \N__37076\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_4_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28781\,
            in1 => \N__26690\,
            in2 => \N__24596\,
            in3 => \N__28091\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_4_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__28440\,
            in1 => \_gnd_net_\,
            in2 => \N__24593\,
            in3 => \N__24467\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_6_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37077\,
            in1 => \_gnd_net_\,
            in2 => \N__24571\,
            in3 => \N__24547\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_4_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__24517\,
            in1 => \N__28778\,
            in2 => \N__26074\,
            in3 => \N__37075\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_4_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28779\,
            in1 => \N__24500\,
            in2 => \N__24485\,
            in3 => \N__24478\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_6_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__28441\,
            in1 => \N__24845\,
            in2 => \N__28974\,
            in3 => \N__24461\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNINA181_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__27749\,
            in1 => \N__31384\,
            in2 => \N__30843\,
            in3 => \N__27988\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27748\,
            in2 => \N__27989\,
            in3 => \N__37089\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__28425\,
            in1 => \N__24680\,
            in2 => \N__24704\,
            in3 => \N__28774\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__24701\,
            in1 => \N__24674\,
            in2 => \N__24692\,
            in3 => \N__28426\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28159\,
            in1 => \_gnd_net_\,
            in2 => \N__37245\,
            in3 => \N__26458\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24667\,
            in1 => \N__26089\,
            in2 => \_gnd_net_\,
            in3 => \N__37088\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIVAI91_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__26090\,
            in1 => \N__31385\,
            in2 => \N__30844\,
            in3 => \N__24668\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI2KHQ1_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__31386\,
            in1 => \N__24656\,
            in2 => \N__24641\,
            in3 => \N__24638\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNI2KHQ1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIPG541_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__24718\,
            in1 => \N__31279\,
            in2 => \N__24836\,
            in3 => \N__30693\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI86UU1_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31280\,
            in1 => \N__24808\,
            in2 => \N__24794\,
            in3 => \N__27002\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI86UU1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQMSM4_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__27251\,
            in2 => \N__24791\,
            in3 => \N__24740\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFG9I8_0_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__27252\,
            in1 => \N__24788\,
            in2 => \N__24782\,
            in3 => \N__24725\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFG9I8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIFAG61_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__30557\,
            in1 => \N__31277\,
            in2 => \N__32651\,
            in3 => \N__30692\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIKPJ32_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31278\,
            in1 => \N__24764\,
            in2 => \N__24743\,
            in3 => \N__31805\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIKPJ32_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI4QLM1_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__26462\,
            in1 => \N__28163\,
            in2 => \N__31536\,
            in3 => \N__24734\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI4QLM1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34907\,
            in1 => \N__32349\,
            in2 => \N__32119\,
            in3 => \N__35988\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33656\,
            ce => \N__24916\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35985\,
            in1 => \N__34911\,
            in2 => \N__39619\,
            in3 => \N__39258\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33656\,
            ce => \N__24916\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34908\,
            in1 => \N__38550\,
            in2 => \N__36194\,
            in3 => \N__38867\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33656\,
            ce => \N__24916\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35986\,
            in1 => \N__34912\,
            in2 => \N__38172\,
            in3 => \N__37755\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33656\,
            ce => \N__24916\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34909\,
            in1 => \N__35189\,
            in2 => \N__36195\,
            in3 => \N__35414\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33656\,
            ce => \N__24916\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__5_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35987\,
            in1 => \N__34913\,
            in2 => \N__30498\,
            in3 => \N__30068\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33656\,
            ce => \N__24916\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34910\,
            in1 => \N__29356\,
            in2 => \N__29643\,
            in3 => \N__35989\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33656\,
            ce => \N__24916\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_6_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37286\,
            in1 => \N__24877\,
            in2 => \_gnd_net_\,
            in3 => \N__24862\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34653\,
            in1 => \N__32399\,
            in2 => \N__32111\,
            in3 => \N__36548\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33665\,
            ce => \N__25087\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36544\,
            in1 => \N__34654\,
            in2 => \N__39636\,
            in3 => \N__39188\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33665\,
            ce => \N__25087\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37411\,
            in1 => \N__26794\,
            in2 => \_gnd_net_\,
            in3 => \N__26812\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__2_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__36545\,
            in1 => \N__38551\,
            in2 => \N__38833\,
            in3 => \N__34657\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33665\,
            ce => \N__25087\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_2_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37410\,
            in1 => \N__26731\,
            in2 => \_gnd_net_\,
            in3 => \N__26752\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36546\,
            in1 => \N__38067\,
            in2 => \N__37857\,
            in3 => \N__34656\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33665\,
            ce => \N__25087\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__4_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36547\,
            in1 => \N__34655\,
            in2 => \N__35548\,
            in3 => \N__35235\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33665\,
            ce => \N__25087\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__26881\,
            in1 => \N__24971\,
            in2 => \N__26861\,
            in3 => \N__28937\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_5_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37450\,
            in1 => \_gnd_net_\,
            in2 => \N__25055\,
            in3 => \N__25034\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_5_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__28561\,
            in1 => \N__26102\,
            in2 => \N__25013\,
            in3 => \N__28939\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_5_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__25010\,
            in1 => \N__24995\,
            in2 => \N__24989\,
            in3 => \N__28562\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26536\,
            in1 => \N__28934\,
            in2 => \N__26519\,
            in3 => \N__37448\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__28938\,
            in1 => \N__24965\,
            in2 => \N__26945\,
            in3 => \N__28560\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25423\,
            in1 => \N__28935\,
            in2 => \N__25406\,
            in3 => \N__37449\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28936\,
            in1 => \N__25390\,
            in2 => \N__25373\,
            in3 => \N__25369\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__4_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34699\,
            in1 => \N__35190\,
            in2 => \N__36599\,
            in3 => \N__35522\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33684\,
            ce => \N__25334\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_4_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__28940\,
            in1 => \N__25129\,
            in2 => \N__25148\,
            in3 => \N__37249\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_4_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26185\,
            in1 => \N__25282\,
            in2 => \N__25262\,
            in3 => \N__28941\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_4_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__28942\,
            in1 => \N__25252\,
            in2 => \N__25237\,
            in3 => \N__37250\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__25216\,
            in1 => \N__25195\,
            in2 => \N__25172\,
            in3 => \N__28943\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_4_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25169\,
            in2 => \N__25163\,
            in3 => \N__28639\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIJRTE1_4_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__31552\,
            in1 => \N__25147\,
            in2 => \N__25133\,
            in3 => \N__30916\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__28637\,
            in1 => \N__25838\,
            in2 => \N__25829\,
            in3 => \N__25472\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__25658\,
            in1 => \N__25814\,
            in2 => \N__25799\,
            in3 => \N__25773\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26342\,
            in1 => \N__25454\,
            in2 => \N__25673\,
            in3 => \N__25659\,
            lcout => \processor_zipi8.sy_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37409\,
            in1 => \N__25504\,
            in2 => \_gnd_net_\,
            in3 => \N__25493\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_2_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__25991\,
            in1 => \N__28633\,
            in2 => \N__25475\,
            in3 => \N__28944\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__28945\,
            in1 => \N__26903\,
            in2 => \N__28657\,
            in3 => \N__25466\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_2_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__38204\,
            in1 => \N__32558\,
            in2 => \N__25457\,
            in3 => \N__28638\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34805\,
            in1 => \N__35885\,
            in2 => \N__32363\,
            in3 => \N__31959\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33702\,
            ce => \N__25957\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000001100"
        )
    port map (
            in0 => \N__39241\,
            in1 => \N__39626\,
            in2 => \N__36098\,
            in3 => \N__34808\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33702\,
            ce => \N__25957\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__34806\,
            in1 => \N__38782\,
            in2 => \N__36099\,
            in3 => \N__38425\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33702\,
            ce => \N__25957\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_2_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25849\,
            in1 => \N__26002\,
            in2 => \_gnd_net_\,
            in3 => \N__37478\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__3_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34807\,
            in1 => \N__35886\,
            in2 => \N__38173\,
            in3 => \N__37629\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33702\,
            ce => \N__25957\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_3_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26200\,
            in1 => \N__25981\,
            in2 => \_gnd_net_\,
            in3 => \N__37477\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__5_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__35884\,
            in1 => \N__30494\,
            in2 => \N__30150\,
            in3 => \N__34809\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33702\,
            ce => \N__25957\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__33926\,
            in1 => \N__36312\,
            in2 => \N__32364\,
            in3 => \N__32058\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33705\,
            ce => \N__26168\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36309\,
            in1 => \N__33929\,
            in2 => \N__39645\,
            in3 => \N__39226\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33705\,
            ce => \N__26168\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__33927\,
            in1 => \N__36313\,
            in2 => \N__38531\,
            in3 => \N__38783\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33705\,
            ce => \N__26168\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36310\,
            in1 => \N__33930\,
            in2 => \N__38186\,
            in3 => \N__37705\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33705\,
            ce => \N__26168\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__33928\,
            in1 => \N__35220\,
            in2 => \N__35568\,
            in3 => \N__36314\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33705\,
            ce => \N__26168\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__5_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36311\,
            in1 => \N__33931\,
            in2 => \N__30510\,
            in3 => \N__30117\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33705\,
            ce => \N__26168\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_5_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26125\,
            in1 => \N__26113\,
            in2 => \_gnd_net_\,
            in3 => \N__37490\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34610\,
            in1 => \N__36619\,
            in2 => \N__32352\,
            in3 => \N__32123\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__1_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36615\,
            in1 => \N__39637\,
            in2 => \N__39284\,
            in3 => \N__34616\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34611\,
            in1 => \N__36620\,
            in2 => \N__38576\,
            in3 => \N__38889\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__3_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36616\,
            in1 => \N__34614\,
            in2 => \N__38192\,
            in3 => \N__37778\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__4_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34612\,
            in1 => \N__36621\,
            in2 => \N__35232\,
            in3 => \N__35428\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__5_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36617\,
            in1 => \N__34615\,
            in2 => \N__30473\,
            in3 => \N__30154\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__6_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34613\,
            in1 => \N__36622\,
            in2 => \N__29368\,
            in3 => \N__29772\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__7_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36618\,
            in1 => \N__33334\,
            in2 => \N__33001\,
            in3 => \N__34617\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33697\,
            ce => \N__26294\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNITG181_3_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__28070\,
            in1 => \N__31515\,
            in2 => \N__30979\,
            in3 => \N__27941\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_3_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37071\,
            in1 => \N__27094\,
            in2 => \_gnd_net_\,
            in3 => \N__28108\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26246\,
            in1 => \N__28527\,
            in2 => \N__26282\,
            in3 => \N__28893\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28528\,
            in1 => \N__26279\,
            in2 => \N__26270\,
            in3 => \N__26240\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_3_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28069\,
            in1 => \N__27940\,
            in2 => \_gnd_net_\,
            in3 => \N__37069\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_3_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37070\,
            in1 => \N__26215\,
            in2 => \_gnd_net_\,
            in3 => \N__26233\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI5HI91_3_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26234\,
            in1 => \N__31516\,
            in2 => \N__26219\,
            in3 => \N__30864\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIE0IQ1_3_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31517\,
            in1 => \N__26390\,
            in2 => \N__26372\,
            in3 => \N__26369\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIE0IQ1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_2_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27808\,
            in1 => \N__26602\,
            in2 => \_gnd_net_\,
            in3 => \N__37066\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIRE181_2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__27716\,
            in1 => \N__31507\,
            in2 => \N__30943\,
            in3 => \N__27950\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27949\,
            in1 => \N__27715\,
            in2 => \_gnd_net_\,
            in3 => \N__37068\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_2_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__28767\,
            in1 => \N__26327\,
            in2 => \N__26354\,
            in3 => \N__28427\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_2_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28428\,
            in1 => \N__26351\,
            in2 => \N__26345\,
            in3 => \N__26321\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_2_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37064\,
            in1 => \_gnd_net_\,
            in2 => \N__28129\,
            in3 => \N__26716\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__27727\,
            in1 => \N__28766\,
            in2 => \N__27967\,
            in3 => \N__37065\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_2_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37067\,
            in1 => \N__26620\,
            in2 => \_gnd_net_\,
            in3 => \N__26647\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34582\,
            in1 => \N__36382\,
            in2 => \N__32474\,
            in3 => \N__32088\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36378\,
            in1 => \N__39608\,
            in2 => \N__39289\,
            in3 => \N__34586\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34583\,
            in1 => \N__36383\,
            in2 => \N__38569\,
            in3 => \N__38800\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36379\,
            in1 => \N__38136\,
            in2 => \N__37835\,
            in3 => \N__34587\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34584\,
            in1 => \N__36384\,
            in2 => \N__35236\,
            in3 => \N__35498\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36380\,
            in1 => \N__30477\,
            in2 => \N__30136\,
            in3 => \N__34588\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34585\,
            in1 => \N__36385\,
            in2 => \N__29395\,
            in3 => \N__29708\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36381\,
            in1 => \N__33290\,
            in2 => \N__32999\,
            in3 => \N__34589\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33666\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIVI181_4_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__30659\,
            in1 => \N__28061\,
            in2 => \N__28244\,
            in3 => \N__31341\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIKAMM1_4_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31342\,
            in1 => \N__26689\,
            in2 => \N__26669\,
            in3 => \N__28084\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIKAMM1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIPC181_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__30656\,
            in1 => \N__27734\,
            in2 => \N__27971\,
            in3 => \N__31337\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI8ULM1_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31338\,
            in1 => \N__26579\,
            in2 => \N__26651\,
            in3 => \N__28142\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI3FI91_2_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__30658\,
            in1 => \N__26648\,
            in2 => \N__26624\,
            in3 => \N__31339\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIASHQ1_2_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31340\,
            in1 => \N__27809\,
            in2 => \N__26606\,
            in3 => \N__26603\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIASHQ1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__28141\,
            in1 => \N__26578\,
            in2 => \N__26564\,
            in3 => \N__28889\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI1DI91_1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__31336\,
            in1 => \N__26540\,
            in2 => \N__26515\,
            in3 => \N__30657\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI2VSM4_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26780\,
            in1 => \N__27191\,
            in2 => \N__26768\,
            in3 => \N__27540\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV0AI8_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__27192\,
            in1 => \N__26489\,
            in2 => \N__26480\,
            in3 => \N__26825\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI6OHQ1_1_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__26891\,
            in1 => \N__26867\,
            in2 => \N__26860\,
            in3 => \N__31175\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIHCG61_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30635\,
            in1 => \N__32621\,
            in2 => \N__31305\,
            in3 => \N__32605\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIRI541_1_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26819\,
            in1 => \N__31172\,
            in2 => \N__26801\,
            in3 => \N__30636\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNICAUU1_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31173\,
            in1 => \N__26978\,
            in2 => \N__26783\,
            in3 => \N__26960\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIOTJ32_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010101"
        )
    port map (
            in0 => \N__26774\,
            in1 => \N__38924\,
            in2 => \N__38948\,
            in3 => \N__31174\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIJEG61_2_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__32570\,
            in1 => \N__31217\,
            in2 => \N__32585\,
            in3 => \N__30690\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIS1K32_2_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__31219\,
            in1 => \N__38219\,
            in2 => \N__26759\,
            in3 => \N__38240\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIS1K32_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNITK541_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26756\,
            in1 => \N__31218\,
            in2 => \N__26741\,
            in3 => \N__30691\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIC2MM1_2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31221\,
            in1 => \N__26720\,
            in2 => \N__26705\,
            in3 => \N__28133\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIC2MM1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFHAI8_2_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__27059\,
            in1 => \N__27008\,
            in2 => \N__27044\,
            in3 => \N__27206\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFHAI8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIGEUU1_2_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31220\,
            in1 => \N__26933\,
            in2 => \N__27026\,
            in3 => \N__26915\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIGEUU1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA7TM4_2_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__27541\,
            in1 => \N__27017\,
            in2 => \N__27011\,
            in3 => \N__27205\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34203\,
            in1 => \N__36185\,
            in2 => \N__32476\,
            in3 => \N__32102\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33686\,
            ce => \N__27686\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36181\,
            in1 => \N__34204\,
            in2 => \N__39542\,
            in3 => \N__39261\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33686\,
            ce => \N__27686\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26977\,
            in1 => \N__26956\,
            in2 => \_gnd_net_\,
            in3 => \N__37432\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__2_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36182\,
            in1 => \N__38831\,
            in2 => \N__38570\,
            in3 => \N__34207\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33686\,
            ce => \N__27686\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_2_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26932\,
            in1 => \N__26914\,
            in2 => \_gnd_net_\,
            in3 => \N__37430\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__3_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36183\,
            in1 => \N__34205\,
            in2 => \N__38182\,
            in3 => \N__37702\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33686\,
            ce => \N__27686\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_3_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27928\,
            in1 => \N__27907\,
            in2 => \_gnd_net_\,
            in3 => \N__37431\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__4_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36184\,
            in1 => \N__34206\,
            in2 => \N__35559\,
            in3 => \N__35170\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33686\,
            ce => \N__27686\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNILGG61_3_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30798\,
            in1 => \N__30536\,
            in2 => \N__31508\,
            in3 => \N__32545\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI06K32_3_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__37538\,
            in1 => \N__37517\,
            in2 => \N__27647\,
            in3 => \N__31326\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI06K32_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIFTM4_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__27896\,
            in1 => \N__27186\,
            in2 => \N__27644\,
            in3 => \N__27539\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV1BI8_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__27187\,
            in1 => \N__27122\,
            in2 => \N__27113\,
            in3 => \N__27065\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV1BI8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIG6MM1_3_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31325\,
            in1 => \N__27095\,
            in2 => \N__27077\,
            in3 => \N__28112\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIG6MM1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIVM541_3_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__27866\,
            in1 => \N__31320\,
            in2 => \N__27890\,
            in3 => \N__30797\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIKIUU1_3_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31321\,
            in1 => \N__27932\,
            in2 => \N__27911\,
            in3 => \N__27908\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIKIUU1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_3_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37438\,
            in2 => \N__32546\,
            in3 => \N__30535\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_3_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27886\,
            in1 => \N__37439\,
            in2 => \_gnd_net_\,
            in3 => \N__27865\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_3_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__27842\,
            in1 => \N__28613\,
            in2 => \N__27833\,
            in3 => \N__28969\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_3_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28614\,
            in1 => \N__36866\,
            in2 => \N__27830\,
            in3 => \N__27827\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__2_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__34726\,
            in1 => \N__38505\,
            in2 => \N__36100\,
            in3 => \N__38832\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33710\,
            ce => \N__27788\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__32120\,
            in1 => \N__32438\,
            in2 => \N__34794\,
            in3 => \N__36847\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36840\,
            in1 => \N__34600\,
            in2 => \N__39646\,
            in3 => \N__39263\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__38882\,
            in1 => \N__36844\,
            in2 => \N__34793\,
            in3 => \N__38574\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__3_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36841\,
            in1 => \N__34601\,
            in2 => \N__38191\,
            in3 => \N__37810\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34598\,
            in1 => \N__36845\,
            in2 => \N__35169\,
            in3 => \N__35545\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36842\,
            in1 => \N__34602\,
            in2 => \N__30514\,
            in3 => \N__30147\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34599\,
            in1 => \N__36846\,
            in2 => \N__29437\,
            in3 => \N__29751\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36843\,
            in1 => \N__33333\,
            in2 => \N__32960\,
            in3 => \N__34609\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33699\,
            ce => \N__28004\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34590\,
            in1 => \N__36740\,
            in2 => \N__32475\,
            in3 => \N__32122\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36736\,
            in1 => \N__34594\,
            in2 => \N__39638\,
            in3 => \N__39243\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34591\,
            in1 => \N__36741\,
            in2 => \N__38888\,
            in3 => \N__38575\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__3_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36737\,
            in1 => \N__34595\,
            in2 => \N__38190\,
            in3 => \N__37756\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34592\,
            in1 => \N__36742\,
            in2 => \N__35233\,
            in3 => \N__35485\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__5_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36738\,
            in1 => \N__34596\,
            in2 => \N__30518\,
            in3 => \N__30148\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__6_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__34593\,
            in1 => \N__36743\,
            in2 => \N__29394\,
            in3 => \N__29710\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__7_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36739\,
            in1 => \N__34597\,
            in2 => \N__33336\,
            in3 => \N__32944\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33688\,
            ce => \N__28181\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__34884\,
            in1 => \N__32461\,
            in2 => \N__36851\,
            in3 => \N__32087\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34885\,
            in1 => \N__39609\,
            in2 => \N__39285\,
            in3 => \N__36830\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__2_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__38541\,
            in1 => \N__34890\,
            in2 => \N__36852\,
            in3 => \N__38801\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__3_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34886\,
            in1 => \N__36819\,
            in2 => \N__38181\,
            in3 => \N__37823\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__4_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__36818\,
            in1 => \N__35221\,
            in2 => \N__35558\,
            in3 => \N__34891\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__5_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__34887\,
            in1 => \N__30481\,
            in2 => \N__30135\,
            in3 => \N__36829\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__6_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__29398\,
            in1 => \N__34889\,
            in2 => \N__36853\,
            in3 => \N__29709\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__7_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__34888\,
            in1 => \N__32872\,
            in2 => \N__33317\,
            in3 => \N__36831\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33677\,
            ce => \N__29036\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_7_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31039\,
            in1 => \N__31060\,
            in2 => \_gnd_net_\,
            in3 => \N__37252\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_7_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37253\,
            in1 => \N__28291\,
            in2 => \_gnd_net_\,
            in3 => \N__28273\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_7_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__31757\,
            in1 => \N__28615\,
            in2 => \N__29018\,
            in3 => \N__29003\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_7_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28616\,
            in1 => \N__28331\,
            in2 => \N__28319\,
            in3 => \N__28316\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI5P181_7_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__30860\,
            in1 => \N__28292\,
            in2 => \N__28277\,
            in3 => \N__31691\,
            lcout => OPEN,
            ltout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI0NMM1_7_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31692\,
            in1 => \N__31768\,
            in2 => \N__28262\,
            in3 => \N__31778\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI0NMM1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_7_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31777\,
            in1 => \_gnd_net_\,
            in2 => \N__31769\,
            in3 => \N__37251\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIDPI91_7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__31690\,
            in1 => \N__31061\,
            in2 => \N__31043\,
            in3 => \N__30859\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34832\,
            in1 => \N__35994\,
            in2 => \N__32458\,
            in3 => \N__32110\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33678\,
            ce => \N__32684\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35990\,
            in1 => \N__34835\,
            in2 => \N__39642\,
            in3 => \N__39177\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33678\,
            ce => \N__32684\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__34833\,
            in1 => \N__38887\,
            in2 => \N__36854\,
            in3 => \N__38565\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33678\,
            ce => \N__32684\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__35991\,
            in1 => \N__38137\,
            in2 => \N__37840\,
            in3 => \N__34838\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33678\,
            ce => \N__32684\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35992\,
            in1 => \N__34836\,
            in2 => \N__30507\,
            in3 => \N__30149\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33678\,
            ce => \N__32684\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34834\,
            in1 => \N__35995\,
            in2 => \N__29768\,
            in3 => \N__29438\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33678\,
            ce => \N__32684\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__7_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__35993\,
            in1 => \N__34837\,
            in2 => \N__33337\,
            in3 => \N__33000\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33678\,
            ce => \N__32684\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34701\,
            in1 => \N__36836\,
            in2 => \N__32459\,
            in3 => \N__32115\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33687\,
            ce => \N__32507\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36832\,
            in1 => \N__34702\,
            in2 => \N__39647\,
            in3 => \N__39242\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33687\,
            ce => \N__32507\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32620\,
            in1 => \N__32606\,
            in2 => \_gnd_net_\,
            in3 => \N__37397\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__2_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36833\,
            in1 => \N__34703\,
            in2 => \N__38843\,
            in3 => \N__38566\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33687\,
            ce => \N__32507\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_2_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32581\,
            in1 => \N__32569\,
            in2 => \_gnd_net_\,
            in3 => \N__37396\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__3_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36834\,
            in1 => \N__38122\,
            in2 => \N__37858\,
            in3 => \N__34831\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33687\,
            ce => \N__32507\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__4_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36835\,
            in1 => \N__34704\,
            in2 => \N__35557\,
            in3 => \N__35240\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33687\,
            ce => \N__32507\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__34198\,
            in1 => \N__36604\,
            in2 => \N__32477\,
            in3 => \N__32101\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33698\,
            ce => \N__33389\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36600\,
            in1 => \N__34199\,
            in2 => \N__39543\,
            in3 => \N__39259\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33698\,
            ce => \N__33389\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38941\,
            in1 => \N__38920\,
            in2 => \_gnd_net_\,
            in3 => \N__37502\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__2_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36601\,
            in1 => \N__34200\,
            in2 => \N__38890\,
            in3 => \N__38549\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33698\,
            ce => \N__33389\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_2_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38236\,
            in1 => \N__38215\,
            in2 => \_gnd_net_\,
            in3 => \N__37500\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__3_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__36602\,
            in1 => \N__34201\,
            in2 => \N__38183\,
            in3 => \N__37836\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33698\,
            ce => \N__33389\,
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_3_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37534\,
            in1 => \N__37516\,
            in2 => \_gnd_net_\,
            in3 => \N__37501\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__4_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__36603\,
            in1 => \N__35531\,
            in2 => \N__35219\,
            in3 => \N__34202\,
            lcout => \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33698\,
            ce => \N__33389\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
