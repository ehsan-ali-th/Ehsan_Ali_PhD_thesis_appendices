// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jul 10 2019 22:39:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    LED1,
    CLK_3P3_MHZ,
    BTN1);

    output LED1;
    input CLK_3P3_MHZ;
    input BTN1;

    wire N__39686;
    wire N__39685;
    wire N__39684;
    wire N__39675;
    wire N__39674;
    wire N__39673;
    wire N__39666;
    wire N__39665;
    wire N__39664;
    wire N__39647;
    wire N__39646;
    wire N__39645;
    wire N__39644;
    wire N__39643;
    wire N__39642;
    wire N__39639;
    wire N__39638;
    wire N__39637;
    wire N__39636;
    wire N__39635;
    wire N__39632;
    wire N__39631;
    wire N__39630;
    wire N__39627;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39609;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39598;
    wire N__39597;
    wire N__39596;
    wire N__39595;
    wire N__39594;
    wire N__39593;
    wire N__39592;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39547;
    wire N__39546;
    wire N__39545;
    wire N__39544;
    wire N__39543;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39503;
    wire N__39498;
    wire N__39495;
    wire N__39494;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39478;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39402;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39369;
    wire N__39366;
    wire N__39359;
    wire N__39350;
    wire N__39345;
    wire N__39342;
    wire N__39335;
    wire N__39330;
    wire N__39321;
    wire N__39318;
    wire N__39313;
    wire N__39308;
    wire N__39303;
    wire N__39290;
    wire N__39289;
    wire N__39286;
    wire N__39285;
    wire N__39284;
    wire N__39283;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39263;
    wire N__39262;
    wire N__39261;
    wire N__39260;
    wire N__39259;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39248;
    wire N__39247;
    wire N__39244;
    wire N__39243;
    wire N__39242;
    wire N__39241;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39233;
    wire N__39230;
    wire N__39229;
    wire N__39228;
    wire N__39227;
    wire N__39226;
    wire N__39225;
    wire N__39224;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39202;
    wire N__39199;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39178;
    wire N__39177;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39131;
    wire N__39128;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39074;
    wire N__39071;
    wire N__39068;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39052;
    wire N__39049;
    wire N__39044;
    wire N__39039;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39015;
    wire N__39012;
    wire N__39007;
    wire N__39000;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38982;
    wire N__38977;
    wire N__38970;
    wire N__38961;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38929;
    wire N__38924;
    wire N__38921;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38890;
    wire N__38889;
    wire N__38888;
    wire N__38887;
    wire N__38886;
    wire N__38883;
    wire N__38882;
    wire N__38881;
    wire N__38880;
    wire N__38879;
    wire N__38878;
    wire N__38875;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38851;
    wire N__38848;
    wire N__38847;
    wire N__38844;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38836;
    wire N__38835;
    wire N__38834;
    wire N__38833;
    wire N__38832;
    wire N__38831;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38821;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38806;
    wire N__38803;
    wire N__38802;
    wire N__38801;
    wire N__38800;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38783;
    wire N__38782;
    wire N__38779;
    wire N__38776;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38761;
    wire N__38758;
    wire N__38755;
    wire N__38752;
    wire N__38747;
    wire N__38744;
    wire N__38739;
    wire N__38732;
    wire N__38731;
    wire N__38730;
    wire N__38729;
    wire N__38726;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38711;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38686;
    wire N__38683;
    wire N__38678;
    wire N__38673;
    wire N__38670;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38648;
    wire N__38641;
    wire N__38636;
    wire N__38633;
    wire N__38626;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38604;
    wire N__38599;
    wire N__38596;
    wire N__38585;
    wire N__38576;
    wire N__38575;
    wire N__38574;
    wire N__38571;
    wire N__38570;
    wire N__38569;
    wire N__38568;
    wire N__38567;
    wire N__38566;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38558;
    wire N__38557;
    wire N__38556;
    wire N__38553;
    wire N__38552;
    wire N__38551;
    wire N__38550;
    wire N__38549;
    wire N__38546;
    wire N__38545;
    wire N__38542;
    wire N__38541;
    wire N__38540;
    wire N__38537;
    wire N__38534;
    wire N__38533;
    wire N__38532;
    wire N__38531;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38519;
    wire N__38518;
    wire N__38517;
    wire N__38514;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38506;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38462;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38447;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38429;
    wire N__38426;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38411;
    wire N__38406;
    wire N__38403;
    wire N__38398;
    wire N__38395;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38368;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38341;
    wire N__38334;
    wire N__38325;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38310;
    wire N__38307;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38289;
    wire N__38282;
    wire N__38279;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38259;
    wire N__38256;
    wire N__38249;
    wire N__38240;
    wire N__38237;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38219;
    wire N__38216;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38191;
    wire N__38190;
    wire N__38189;
    wire N__38188;
    wire N__38187;
    wire N__38186;
    wire N__38185;
    wire N__38184;
    wire N__38183;
    wire N__38182;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38174;
    wire N__38173;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38159;
    wire N__38158;
    wire N__38155;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38147;
    wire N__38146;
    wire N__38145;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38137;
    wire N__38136;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38122;
    wire N__38119;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38099;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38079;
    wire N__38078;
    wire N__38075;
    wire N__38072;
    wire N__38071;
    wire N__38068;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37969;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37939;
    wire N__37936;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37910;
    wire N__37903;
    wire N__37900;
    wire N__37899;
    wire N__37890;
    wire N__37881;
    wire N__37874;
    wire N__37871;
    wire N__37862;
    wire N__37859;
    wire N__37858;
    wire N__37857;
    wire N__37854;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37840;
    wire N__37837;
    wire N__37836;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37825;
    wire N__37824;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37810;
    wire N__37807;
    wire N__37802;
    wire N__37801;
    wire N__37798;
    wire N__37797;
    wire N__37794;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37782;
    wire N__37779;
    wire N__37778;
    wire N__37775;
    wire N__37774;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37756;
    wire N__37755;
    wire N__37754;
    wire N__37753;
    wire N__37750;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37727;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37706;
    wire N__37705;
    wire N__37704;
    wire N__37703;
    wire N__37702;
    wire N__37701;
    wire N__37698;
    wire N__37693;
    wire N__37690;
    wire N__37685;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37669;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37661;
    wire N__37658;
    wire N__37655;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37641;
    wire N__37630;
    wire N__37629;
    wire N__37628;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37570;
    wire N__37565;
    wire N__37560;
    wire N__37555;
    wire N__37538;
    wire N__37535;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37516;
    wire N__37513;
    wire N__37510;
    wire N__37505;
    wire N__37504;
    wire N__37503;
    wire N__37502;
    wire N__37501;
    wire N__37500;
    wire N__37499;
    wire N__37498;
    wire N__37497;
    wire N__37496;
    wire N__37495;
    wire N__37494;
    wire N__37491;
    wire N__37490;
    wire N__37489;
    wire N__37488;
    wire N__37487;
    wire N__37486;
    wire N__37485;
    wire N__37484;
    wire N__37479;
    wire N__37478;
    wire N__37477;
    wire N__37470;
    wire N__37469;
    wire N__37468;
    wire N__37467;
    wire N__37462;
    wire N__37457;
    wire N__37452;
    wire N__37451;
    wire N__37450;
    wire N__37449;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37441;
    wire N__37440;
    wire N__37439;
    wire N__37438;
    wire N__37433;
    wire N__37432;
    wire N__37431;
    wire N__37430;
    wire N__37429;
    wire N__37428;
    wire N__37427;
    wire N__37426;
    wire N__37425;
    wire N__37424;
    wire N__37423;
    wire N__37420;
    wire N__37417;
    wire N__37412;
    wire N__37411;
    wire N__37410;
    wire N__37409;
    wire N__37406;
    wire N__37401;
    wire N__37398;
    wire N__37397;
    wire N__37396;
    wire N__37395;
    wire N__37394;
    wire N__37391;
    wire N__37386;
    wire N__37385;
    wire N__37384;
    wire N__37383;
    wire N__37382;
    wire N__37381;
    wire N__37378;
    wire N__37373;
    wire N__37372;
    wire N__37369;
    wire N__37362;
    wire N__37357;
    wire N__37356;
    wire N__37355;
    wire N__37354;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37333;
    wire N__37332;
    wire N__37331;
    wire N__37330;
    wire N__37329;
    wire N__37328;
    wire N__37327;
    wire N__37324;
    wire N__37323;
    wire N__37322;
    wire N__37317;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37303;
    wire N__37302;
    wire N__37301;
    wire N__37300;
    wire N__37299;
    wire N__37298;
    wire N__37297;
    wire N__37296;
    wire N__37295;
    wire N__37294;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37286;
    wire N__37281;
    wire N__37278;
    wire N__37273;
    wire N__37270;
    wire N__37265;
    wire N__37260;
    wire N__37255;
    wire N__37254;
    wire N__37253;
    wire N__37252;
    wire N__37251;
    wire N__37250;
    wire N__37249;
    wire N__37246;
    wire N__37245;
    wire N__37236;
    wire N__37231;
    wire N__37228;
    wire N__37221;
    wire N__37218;
    wire N__37217;
    wire N__37216;
    wire N__37215;
    wire N__37214;
    wire N__37213;
    wire N__37212;
    wire N__37211;
    wire N__37206;
    wire N__37203;
    wire N__37194;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37172;
    wire N__37163;
    wire N__37154;
    wire N__37147;
    wire N__37140;
    wire N__37137;
    wire N__37136;
    wire N__37135;
    wire N__37134;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37118;
    wire N__37113;
    wire N__37108;
    wire N__37105;
    wire N__37098;
    wire N__37093;
    wire N__37090;
    wire N__37089;
    wire N__37088;
    wire N__37085;
    wire N__37084;
    wire N__37083;
    wire N__37082;
    wire N__37081;
    wire N__37080;
    wire N__37079;
    wire N__37078;
    wire N__37077;
    wire N__37076;
    wire N__37075;
    wire N__37072;
    wire N__37071;
    wire N__37070;
    wire N__37069;
    wire N__37068;
    wire N__37067;
    wire N__37066;
    wire N__37065;
    wire N__37064;
    wire N__37061;
    wire N__37054;
    wire N__37049;
    wire N__37044;
    wire N__37037;
    wire N__37034;
    wire N__37029;
    wire N__37012;
    wire N__37009;
    wire N__37002;
    wire N__36991;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36970;
    wire N__36963;
    wire N__36954;
    wire N__36947;
    wire N__36944;
    wire N__36937;
    wire N__36926;
    wire N__36919;
    wire N__36908;
    wire N__36901;
    wire N__36890;
    wire N__36885;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36853;
    wire N__36852;
    wire N__36851;
    wire N__36850;
    wire N__36849;
    wire N__36848;
    wire N__36847;
    wire N__36846;
    wire N__36845;
    wire N__36844;
    wire N__36843;
    wire N__36842;
    wire N__36841;
    wire N__36840;
    wire N__36837;
    wire N__36836;
    wire N__36835;
    wire N__36834;
    wire N__36833;
    wire N__36832;
    wire N__36831;
    wire N__36830;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36819;
    wire N__36818;
    wire N__36815;
    wire N__36814;
    wire N__36813;
    wire N__36812;
    wire N__36811;
    wire N__36810;
    wire N__36809;
    wire N__36808;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36800;
    wire N__36799;
    wire N__36798;
    wire N__36797;
    wire N__36796;
    wire N__36795;
    wire N__36794;
    wire N__36793;
    wire N__36792;
    wire N__36775;
    wire N__36772;
    wire N__36761;
    wire N__36744;
    wire N__36743;
    wire N__36742;
    wire N__36741;
    wire N__36740;
    wire N__36739;
    wire N__36738;
    wire N__36737;
    wire N__36736;
    wire N__36733;
    wire N__36716;
    wire N__36713;
    wire N__36712;
    wire N__36711;
    wire N__36710;
    wire N__36709;
    wire N__36708;
    wire N__36707;
    wire N__36706;
    wire N__36705;
    wire N__36702;
    wire N__36701;
    wire N__36700;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36696;
    wire N__36695;
    wire N__36694;
    wire N__36693;
    wire N__36692;
    wire N__36689;
    wire N__36688;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36668;
    wire N__36667;
    wire N__36666;
    wire N__36665;
    wire N__36664;
    wire N__36663;
    wire N__36662;
    wire N__36661;
    wire N__36660;
    wire N__36659;
    wire N__36658;
    wire N__36657;
    wire N__36656;
    wire N__36655;
    wire N__36652;
    wire N__36645;
    wire N__36628;
    wire N__36627;
    wire N__36626;
    wire N__36625;
    wire N__36624;
    wire N__36623;
    wire N__36622;
    wire N__36621;
    wire N__36620;
    wire N__36619;
    wire N__36618;
    wire N__36617;
    wire N__36616;
    wire N__36615;
    wire N__36614;
    wire N__36613;
    wire N__36612;
    wire N__36611;
    wire N__36610;
    wire N__36609;
    wire N__36608;
    wire N__36607;
    wire N__36606;
    wire N__36605;
    wire N__36604;
    wire N__36603;
    wire N__36602;
    wire N__36601;
    wire N__36600;
    wire N__36599;
    wire N__36598;
    wire N__36597;
    wire N__36596;
    wire N__36595;
    wire N__36594;
    wire N__36593;
    wire N__36588;
    wire N__36585;
    wire N__36568;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36558;
    wire N__36557;
    wire N__36556;
    wire N__36555;
    wire N__36554;
    wire N__36553;
    wire N__36552;
    wire N__36551;
    wire N__36550;
    wire N__36549;
    wire N__36548;
    wire N__36547;
    wire N__36546;
    wire N__36545;
    wire N__36544;
    wire N__36527;
    wire N__36526;
    wire N__36525;
    wire N__36524;
    wire N__36523;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36503;
    wire N__36502;
    wire N__36501;
    wire N__36488;
    wire N__36485;
    wire N__36484;
    wire N__36477;
    wire N__36470;
    wire N__36467;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36455;
    wire N__36450;
    wire N__36447;
    wire N__36430;
    wire N__36415;
    wire N__36414;
    wire N__36413;
    wire N__36412;
    wire N__36411;
    wire N__36410;
    wire N__36407;
    wire N__36406;
    wire N__36405;
    wire N__36404;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36386;
    wire N__36385;
    wire N__36384;
    wire N__36383;
    wire N__36382;
    wire N__36381;
    wire N__36380;
    wire N__36379;
    wire N__36378;
    wire N__36377;
    wire N__36374;
    wire N__36373;
    wire N__36372;
    wire N__36371;
    wire N__36370;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36366;
    wire N__36353;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36333;
    wire N__36316;
    wire N__36315;
    wire N__36314;
    wire N__36313;
    wire N__36312;
    wire N__36311;
    wire N__36310;
    wire N__36309;
    wire N__36298;
    wire N__36295;
    wire N__36288;
    wire N__36285;
    wire N__36284;
    wire N__36283;
    wire N__36282;
    wire N__36281;
    wire N__36280;
    wire N__36279;
    wire N__36276;
    wire N__36263;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36223;
    wire N__36218;
    wire N__36207;
    wire N__36204;
    wire N__36203;
    wire N__36202;
    wire N__36201;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36191;
    wire N__36190;
    wire N__36189;
    wire N__36188;
    wire N__36187;
    wire N__36186;
    wire N__36185;
    wire N__36184;
    wire N__36183;
    wire N__36182;
    wire N__36181;
    wire N__36168;
    wire N__36165;
    wire N__36148;
    wire N__36145;
    wire N__36144;
    wire N__36143;
    wire N__36142;
    wire N__36141;
    wire N__36140;
    wire N__36139;
    wire N__36138;
    wire N__36137;
    wire N__36134;
    wire N__36117;
    wire N__36112;
    wire N__36103;
    wire N__36102;
    wire N__36101;
    wire N__36100;
    wire N__36099;
    wire N__36098;
    wire N__36095;
    wire N__36082;
    wire N__36079;
    wire N__36074;
    wire N__36071;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36051;
    wire N__36050;
    wire N__36035;
    wire N__36034;
    wire N__36029;
    wire N__36024;
    wire N__36019;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35995;
    wire N__35994;
    wire N__35993;
    wire N__35992;
    wire N__35991;
    wire N__35990;
    wire N__35989;
    wire N__35988;
    wire N__35987;
    wire N__35986;
    wire N__35985;
    wire N__35984;
    wire N__35983;
    wire N__35982;
    wire N__35981;
    wire N__35980;
    wire N__35979;
    wire N__35978;
    wire N__35977;
    wire N__35976;
    wire N__35975;
    wire N__35974;
    wire N__35973;
    wire N__35972;
    wire N__35971;
    wire N__35970;
    wire N__35969;
    wire N__35952;
    wire N__35941;
    wire N__35934;
    wire N__35931;
    wire N__35926;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35887;
    wire N__35886;
    wire N__35885;
    wire N__35884;
    wire N__35883;
    wire N__35882;
    wire N__35881;
    wire N__35880;
    wire N__35879;
    wire N__35878;
    wire N__35877;
    wire N__35876;
    wire N__35871;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35854;
    wire N__35849;
    wire N__35848;
    wire N__35847;
    wire N__35846;
    wire N__35845;
    wire N__35844;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35832;
    wire N__35827;
    wire N__35822;
    wire N__35809;
    wire N__35798;
    wire N__35791;
    wire N__35778;
    wire N__35763;
    wire N__35758;
    wire N__35755;
    wire N__35750;
    wire N__35747;
    wire N__35746;
    wire N__35745;
    wire N__35742;
    wire N__35737;
    wire N__35732;
    wire N__35731;
    wire N__35730;
    wire N__35727;
    wire N__35724;
    wire N__35715;
    wire N__35698;
    wire N__35693;
    wire N__35686;
    wire N__35681;
    wire N__35668;
    wire N__35663;
    wire N__35658;
    wire N__35649;
    wire N__35644;
    wire N__35637;
    wire N__35634;
    wire N__35629;
    wire N__35622;
    wire N__35617;
    wire N__35600;
    wire N__35593;
    wire N__35588;
    wire N__35573;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35560;
    wire N__35559;
    wire N__35558;
    wire N__35557;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35549;
    wire N__35548;
    wire N__35547;
    wire N__35546;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35535;
    wire N__35532;
    wire N__35531;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35523;
    wire N__35522;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35498;
    wire N__35495;
    wire N__35494;
    wire N__35489;
    wire N__35486;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35423;
    wire N__35418;
    wire N__35415;
    wire N__35414;
    wire N__35413;
    wire N__35410;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35382;
    wire N__35377;
    wire N__35372;
    wire N__35367;
    wire N__35364;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35340;
    wire N__35333;
    wire N__35328;
    wire N__35319;
    wire N__35314;
    wire N__35311;
    wire N__35306;
    wire N__35303;
    wire N__35298;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35280;
    wire N__35275;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35255;
    wire N__35240;
    wire N__35237;
    wire N__35236;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35231;
    wire N__35230;
    wire N__35229;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35221;
    wire N__35220;
    wire N__35219;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35204;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35193;
    wire N__35192;
    wire N__35191;
    wire N__35190;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35171;
    wire N__35170;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35156;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35123;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35090;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35032;
    wire N__35029;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35008;
    wire N__35007;
    wire N__35006;
    wire N__35001;
    wire N__34996;
    wire N__34989;
    wire N__34986;
    wire N__34979;
    wire N__34968;
    wire N__34965;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34940;
    wire N__34935;
    wire N__34926;
    wire N__34913;
    wire N__34912;
    wire N__34911;
    wire N__34910;
    wire N__34909;
    wire N__34908;
    wire N__34907;
    wire N__34892;
    wire N__34891;
    wire N__34890;
    wire N__34889;
    wire N__34888;
    wire N__34887;
    wire N__34886;
    wire N__34885;
    wire N__34884;
    wire N__34883;
    wire N__34882;
    wire N__34881;
    wire N__34880;
    wire N__34877;
    wire N__34862;
    wire N__34859;
    wire N__34852;
    wire N__34851;
    wire N__34850;
    wire N__34847;
    wire N__34846;
    wire N__34845;
    wire N__34844;
    wire N__34843;
    wire N__34842;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34838;
    wire N__34837;
    wire N__34836;
    wire N__34835;
    wire N__34834;
    wire N__34833;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34829;
    wire N__34828;
    wire N__34827;
    wire N__34826;
    wire N__34825;
    wire N__34824;
    wire N__34823;
    wire N__34822;
    wire N__34821;
    wire N__34820;
    wire N__34819;
    wire N__34818;
    wire N__34817;
    wire N__34816;
    wire N__34815;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34811;
    wire N__34810;
    wire N__34809;
    wire N__34808;
    wire N__34807;
    wire N__34806;
    wire N__34805;
    wire N__34804;
    wire N__34803;
    wire N__34802;
    wire N__34801;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34794;
    wire N__34793;
    wire N__34786;
    wire N__34783;
    wire N__34766;
    wire N__34765;
    wire N__34764;
    wire N__34761;
    wire N__34760;
    wire N__34757;
    wire N__34756;
    wire N__34755;
    wire N__34754;
    wire N__34753;
    wire N__34752;
    wire N__34751;
    wire N__34748;
    wire N__34747;
    wire N__34746;
    wire N__34745;
    wire N__34744;
    wire N__34743;
    wire N__34742;
    wire N__34727;
    wire N__34726;
    wire N__34723;
    wire N__34712;
    wire N__34711;
    wire N__34708;
    wire N__34705;
    wire N__34704;
    wire N__34703;
    wire N__34702;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34686;
    wire N__34669;
    wire N__34658;
    wire N__34657;
    wire N__34656;
    wire N__34655;
    wire N__34654;
    wire N__34653;
    wire N__34640;
    wire N__34639;
    wire N__34638;
    wire N__34637;
    wire N__34636;
    wire N__34635;
    wire N__34634;
    wire N__34633;
    wire N__34626;
    wire N__34625;
    wire N__34624;
    wire N__34621;
    wire N__34620;
    wire N__34619;
    wire N__34618;
    wire N__34617;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34602;
    wire N__34601;
    wire N__34600;
    wire N__34599;
    wire N__34598;
    wire N__34597;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34592;
    wire N__34591;
    wire N__34590;
    wire N__34589;
    wire N__34588;
    wire N__34587;
    wire N__34586;
    wire N__34585;
    wire N__34584;
    wire N__34583;
    wire N__34582;
    wire N__34581;
    wire N__34580;
    wire N__34579;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34553;
    wire N__34536;
    wire N__34521;
    wire N__34520;
    wire N__34519;
    wire N__34518;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34505;
    wire N__34504;
    wire N__34503;
    wire N__34502;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34496;
    wire N__34495;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34478;
    wire N__34469;
    wire N__34468;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34454;
    wire N__34443;
    wire N__34440;
    wire N__34425;
    wire N__34422;
    wire N__34409;
    wire N__34408;
    wire N__34407;
    wire N__34406;
    wire N__34405;
    wire N__34404;
    wire N__34403;
    wire N__34402;
    wire N__34385;
    wire N__34368;
    wire N__34351;
    wire N__34334;
    wire N__34327;
    wire N__34326;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34307;
    wire N__34306;
    wire N__34305;
    wire N__34304;
    wire N__34303;
    wire N__34300;
    wire N__34287;
    wire N__34280;
    wire N__34277;
    wire N__34276;
    wire N__34267;
    wire N__34264;
    wire N__34247;
    wire N__34230;
    wire N__34227;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34211;
    wire N__34208;
    wire N__34207;
    wire N__34206;
    wire N__34205;
    wire N__34204;
    wire N__34203;
    wire N__34202;
    wire N__34201;
    wire N__34200;
    wire N__34199;
    wire N__34198;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34190;
    wire N__34189;
    wire N__34188;
    wire N__34187;
    wire N__34184;
    wire N__34183;
    wire N__34182;
    wire N__34181;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34167;
    wire N__34158;
    wire N__34143;
    wire N__34134;
    wire N__34131;
    wire N__34130;
    wire N__34129;
    wire N__34128;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34097;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34085;
    wire N__34084;
    wire N__34083;
    wire N__34082;
    wire N__34081;
    wire N__34080;
    wire N__34079;
    wire N__34078;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34072;
    wire N__34071;
    wire N__34070;
    wire N__34069;
    wire N__34068;
    wire N__34059;
    wire N__34054;
    wire N__34045;
    wire N__34034;
    wire N__34023;
    wire N__34006;
    wire N__34003;
    wire N__33988;
    wire N__33979;
    wire N__33976;
    wire N__33971;
    wire N__33968;
    wire N__33963;
    wire N__33960;
    wire N__33955;
    wire N__33954;
    wire N__33953;
    wire N__33952;
    wire N__33951;
    wire N__33950;
    wire N__33949;
    wire N__33948;
    wire N__33947;
    wire N__33932;
    wire N__33931;
    wire N__33930;
    wire N__33929;
    wire N__33928;
    wire N__33927;
    wire N__33926;
    wire N__33921;
    wire N__33914;
    wire N__33909;
    wire N__33908;
    wire N__33905;
    wire N__33904;
    wire N__33903;
    wire N__33902;
    wire N__33899;
    wire N__33884;
    wire N__33879;
    wire N__33870;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33858;
    wire N__33855;
    wire N__33846;
    wire N__33829;
    wire N__33826;
    wire N__33825;
    wire N__33824;
    wire N__33823;
    wire N__33810;
    wire N__33803;
    wire N__33792;
    wire N__33787;
    wire N__33782;
    wire N__33779;
    wire N__33772;
    wire N__33763;
    wire N__33760;
    wire N__33755;
    wire N__33750;
    wire N__33731;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33709;
    wire N__33708;
    wire N__33707;
    wire N__33706;
    wire N__33705;
    wire N__33704;
    wire N__33703;
    wire N__33702;
    wire N__33701;
    wire N__33700;
    wire N__33699;
    wire N__33698;
    wire N__33697;
    wire N__33696;
    wire N__33695;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33691;
    wire N__33690;
    wire N__33689;
    wire N__33688;
    wire N__33687;
    wire N__33686;
    wire N__33685;
    wire N__33684;
    wire N__33683;
    wire N__33682;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33677;
    wire N__33676;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33669;
    wire N__33668;
    wire N__33667;
    wire N__33666;
    wire N__33665;
    wire N__33664;
    wire N__33663;
    wire N__33662;
    wire N__33661;
    wire N__33660;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33655;
    wire N__33654;
    wire N__33653;
    wire N__33652;
    wire N__33651;
    wire N__33650;
    wire N__33649;
    wire N__33648;
    wire N__33647;
    wire N__33646;
    wire N__33645;
    wire N__33644;
    wire N__33643;
    wire N__33642;
    wire N__33641;
    wire N__33640;
    wire N__33639;
    wire N__33638;
    wire N__33637;
    wire N__33636;
    wire N__33635;
    wire N__33634;
    wire N__33633;
    wire N__33632;
    wire N__33631;
    wire N__33630;
    wire N__33629;
    wire N__33628;
    wire N__33627;
    wire N__33626;
    wire N__33625;
    wire N__33624;
    wire N__33623;
    wire N__33622;
    wire N__33621;
    wire N__33620;
    wire N__33619;
    wire N__33618;
    wire N__33617;
    wire N__33616;
    wire N__33615;
    wire N__33614;
    wire N__33613;
    wire N__33612;
    wire N__33611;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33606;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33359;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33342;
    wire N__33341;
    wire N__33340;
    wire N__33339;
    wire N__33338;
    wire N__33337;
    wire N__33336;
    wire N__33335;
    wire N__33334;
    wire N__33333;
    wire N__33328;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33317;
    wire N__33316;
    wire N__33313;
    wire N__33312;
    wire N__33311;
    wire N__33310;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33302;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33294;
    wire N__33291;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33267;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33203;
    wire N__33194;
    wire N__33191;
    wire N__33186;
    wire N__33183;
    wire N__33178;
    wire N__33175;
    wire N__33174;
    wire N__33171;
    wire N__33164;
    wire N__33161;
    wire N__33148;
    wire N__33147;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33080;
    wire N__33077;
    wire N__33072;
    wire N__33067;
    wire N__33062;
    wire N__33059;
    wire N__33054;
    wire N__33051;
    wire N__33040;
    wire N__33029;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33021;
    wire N__33018;
    wire N__33017;
    wire N__33016;
    wire N__33015;
    wire N__33014;
    wire N__33013;
    wire N__33012;
    wire N__33011;
    wire N__33010;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33002;
    wire N__33001;
    wire N__33000;
    wire N__32999;
    wire N__32996;
    wire N__32995;
    wire N__32994;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32980;
    wire N__32979;
    wire N__32978;
    wire N__32975;
    wire N__32974;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32876;
    wire N__32873;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32849;
    wire N__32838;
    wire N__32835;
    wire N__32828;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32812;
    wire N__32809;
    wire N__32804;
    wire N__32801;
    wire N__32794;
    wire N__32793;
    wire N__32792;
    wire N__32777;
    wire N__32772;
    wire N__32769;
    wire N__32762;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32741;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32723;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32668;
    wire N__32665;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32651;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32621;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32606;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32581;
    wire N__32578;
    wire N__32575;
    wire N__32570;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32524;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32477;
    wire N__32476;
    wire N__32475;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32455;
    wire N__32452;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32439;
    wire N__32438;
    wire N__32437;
    wire N__32434;
    wire N__32433;
    wire N__32432;
    wire N__32431;
    wire N__32428;
    wire N__32423;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32403;
    wire N__32400;
    wire N__32399;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32381;
    wire N__32380;
    wire N__32377;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32364;
    wire N__32363;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32352;
    wire N__32351;
    wire N__32350;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32335;
    wire N__32332;
    wire N__32325;
    wire N__32324;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32300;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32289;
    wire N__32286;
    wire N__32279;
    wire N__32276;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32264;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32245;
    wire N__32244;
    wire N__32241;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32168;
    wire N__32165;
    wire N__32160;
    wire N__32153;
    wire N__32144;
    wire N__32141;
    wire N__32136;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32120;
    wire N__32119;
    wire N__32116;
    wire N__32115;
    wire N__32112;
    wire N__32111;
    wire N__32110;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32102;
    wire N__32101;
    wire N__32100;
    wire N__32099;
    wire N__32098;
    wire N__32097;
    wire N__32094;
    wire N__32093;
    wire N__32092;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32080;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31997;
    wire N__31992;
    wire N__31989;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31968;
    wire N__31963;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31898;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31871;
    wire N__31868;
    wire N__31863;
    wire N__31858;
    wire N__31851;
    wire N__31842;
    wire N__31841;
    wire N__31832;
    wire N__31827;
    wire N__31824;
    wire N__31819;
    wire N__31816;
    wire N__31805;
    wire N__31802;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31778;
    wire N__31777;
    wire N__31772;
    wire N__31769;
    wire N__31768;
    wire N__31765;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31750;
    wire N__31749;
    wire N__31746;
    wire N__31745;
    wire N__31744;
    wire N__31743;
    wire N__31742;
    wire N__31741;
    wire N__31738;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31734;
    wire N__31733;
    wire N__31732;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31718;
    wire N__31717;
    wire N__31714;
    wire N__31713;
    wire N__31712;
    wire N__31709;
    wire N__31708;
    wire N__31707;
    wire N__31706;
    wire N__31705;
    wire N__31704;
    wire N__31703;
    wire N__31702;
    wire N__31701;
    wire N__31700;
    wire N__31699;
    wire N__31698;
    wire N__31697;
    wire N__31696;
    wire N__31695;
    wire N__31694;
    wire N__31693;
    wire N__31692;
    wire N__31691;
    wire N__31690;
    wire N__31689;
    wire N__31688;
    wire N__31685;
    wire N__31684;
    wire N__31683;
    wire N__31682;
    wire N__31681;
    wire N__31680;
    wire N__31679;
    wire N__31678;
    wire N__31677;
    wire N__31676;
    wire N__31675;
    wire N__31674;
    wire N__31673;
    wire N__31664;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31652;
    wire N__31647;
    wire N__31642;
    wire N__31639;
    wire N__31632;
    wire N__31625;
    wire N__31624;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31616;
    wire N__31615;
    wire N__31614;
    wire N__31613;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31586;
    wire N__31585;
    wire N__31584;
    wire N__31583;
    wire N__31582;
    wire N__31581;
    wire N__31578;
    wire N__31577;
    wire N__31576;
    wire N__31575;
    wire N__31574;
    wire N__31573;
    wire N__31572;
    wire N__31571;
    wire N__31570;
    wire N__31569;
    wire N__31568;
    wire N__31565;
    wire N__31558;
    wire N__31553;
    wire N__31552;
    wire N__31549;
    wire N__31542;
    wire N__31541;
    wire N__31540;
    wire N__31539;
    wire N__31538;
    wire N__31537;
    wire N__31536;
    wire N__31525;
    wire N__31518;
    wire N__31517;
    wire N__31516;
    wire N__31515;
    wire N__31514;
    wire N__31513;
    wire N__31512;
    wire N__31509;
    wire N__31508;
    wire N__31507;
    wire N__31504;
    wire N__31497;
    wire N__31490;
    wire N__31483;
    wire N__31472;
    wire N__31463;
    wire N__31454;
    wire N__31449;
    wire N__31440;
    wire N__31429;
    wire N__31428;
    wire N__31427;
    wire N__31426;
    wire N__31425;
    wire N__31424;
    wire N__31421;
    wire N__31414;
    wire N__31409;
    wire N__31404;
    wire N__31399;
    wire N__31398;
    wire N__31395;
    wire N__31394;
    wire N__31393;
    wire N__31392;
    wire N__31391;
    wire N__31390;
    wire N__31387;
    wire N__31386;
    wire N__31385;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31370;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31343;
    wire N__31342;
    wire N__31341;
    wire N__31340;
    wire N__31339;
    wire N__31338;
    wire N__31337;
    wire N__31336;
    wire N__31327;
    wire N__31326;
    wire N__31325;
    wire N__31322;
    wire N__31321;
    wire N__31320;
    wire N__31317;
    wire N__31306;
    wire N__31305;
    wire N__31302;
    wire N__31297;
    wire N__31292;
    wire N__31281;
    wire N__31280;
    wire N__31279;
    wire N__31278;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31264;
    wire N__31255;
    wire N__31248;
    wire N__31245;
    wire N__31238;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31221;
    wire N__31220;
    wire N__31219;
    wire N__31218;
    wire N__31217;
    wire N__31210;
    wire N__31195;
    wire N__31192;
    wire N__31181;
    wire N__31176;
    wire N__31175;
    wire N__31174;
    wire N__31173;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31159;
    wire N__31150;
    wire N__31141;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31123;
    wire N__31112;
    wire N__31107;
    wire N__31100;
    wire N__31089;
    wire N__31078;
    wire N__31061;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31021;
    wire N__31018;
    wire N__31017;
    wire N__31016;
    wire N__31015;
    wire N__31014;
    wire N__31013;
    wire N__31010;
    wire N__31009;
    wire N__31008;
    wire N__31007;
    wire N__31006;
    wire N__31005;
    wire N__31004;
    wire N__31001;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30986;
    wire N__30985;
    wire N__30984;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30980;
    wire N__30979;
    wire N__30976;
    wire N__30975;
    wire N__30974;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30962;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30946;
    wire N__30945;
    wire N__30944;
    wire N__30943;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30932;
    wire N__30931;
    wire N__30928;
    wire N__30923;
    wire N__30922;
    wire N__30921;
    wire N__30918;
    wire N__30917;
    wire N__30916;
    wire N__30911;
    wire N__30910;
    wire N__30909;
    wire N__30904;
    wire N__30901;
    wire N__30900;
    wire N__30899;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30887;
    wire N__30882;
    wire N__30877;
    wire N__30870;
    wire N__30865;
    wire N__30864;
    wire N__30861;
    wire N__30860;
    wire N__30859;
    wire N__30856;
    wire N__30849;
    wire N__30848;
    wire N__30847;
    wire N__30846;
    wire N__30845;
    wire N__30844;
    wire N__30843;
    wire N__30838;
    wire N__30837;
    wire N__30836;
    wire N__30835;
    wire N__30834;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30823;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30802;
    wire N__30799;
    wire N__30798;
    wire N__30797;
    wire N__30794;
    wire N__30787;
    wire N__30780;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30749;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30730;
    wire N__30723;
    wire N__30716;
    wire N__30709;
    wire N__30704;
    wire N__30699;
    wire N__30694;
    wire N__30693;
    wire N__30692;
    wire N__30691;
    wire N__30690;
    wire N__30685;
    wire N__30682;
    wire N__30675;
    wire N__30670;
    wire N__30667;
    wire N__30660;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30656;
    wire N__30653;
    wire N__30648;
    wire N__30637;
    wire N__30636;
    wire N__30635;
    wire N__30628;
    wire N__30623;
    wire N__30618;
    wire N__30609;
    wire N__30604;
    wire N__30595;
    wire N__30588;
    wire N__30583;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30536;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30514;
    wire N__30511;
    wire N__30510;
    wire N__30509;
    wire N__30508;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30500;
    wire N__30499;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30493;
    wire N__30492;
    wire N__30491;
    wire N__30490;
    wire N__30489;
    wire N__30486;
    wire N__30485;
    wire N__30482;
    wire N__30481;
    wire N__30478;
    wire N__30477;
    wire N__30474;
    wire N__30473;
    wire N__30472;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30464;
    wire N__30463;
    wire N__30462;
    wire N__30461;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30448;
    wire N__30445;
    wire N__30444;
    wire N__30441;
    wire N__30440;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30395;
    wire N__30394;
    wire N__30391;
    wire N__30390;
    wire N__30387;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30288;
    wire N__30281;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30269;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30224;
    wire N__30219;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30207;
    wire N__30204;
    wire N__30197;
    wire N__30192;
    wire N__30187;
    wire N__30178;
    wire N__30173;
    wire N__30170;
    wire N__30155;
    wire N__30154;
    wire N__30151;
    wire N__30150;
    wire N__30149;
    wire N__30148;
    wire N__30147;
    wire N__30146;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30137;
    wire N__30136;
    wire N__30135;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30121;
    wire N__30118;
    wire N__30117;
    wire N__30116;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30090;
    wire N__30089;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30077;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30069;
    wire N__30068;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30057;
    wire N__30048;
    wire N__30045;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30024;
    wire N__30021;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29982;
    wire N__29979;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29952;
    wire N__29951;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29937;
    wire N__29928;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29878;
    wire N__29875;
    wire N__29866;
    wire N__29861;
    wire N__29856;
    wire N__29853;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29834;
    wire N__29831;
    wire N__29816;
    wire N__29813;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29783;
    wire N__29782;
    wire N__29781;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29773;
    wire N__29772;
    wire N__29771;
    wire N__29770;
    wire N__29769;
    wire N__29768;
    wire N__29765;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29744;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29736;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29722;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29710;
    wire N__29709;
    wire N__29708;
    wire N__29707;
    wire N__29706;
    wire N__29705;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29672;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29643;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29633;
    wire N__29630;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29586;
    wire N__29581;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29554;
    wire N__29553;
    wire N__29548;
    wire N__29541;
    wire N__29538;
    wire N__29529;
    wire N__29524;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29485;
    wire N__29480;
    wire N__29477;
    wire N__29470;
    wire N__29467;
    wire N__29460;
    wire N__29447;
    wire N__29446;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29438;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29408;
    wire N__29407;
    wire N__29406;
    wire N__29399;
    wire N__29398;
    wire N__29397;
    wire N__29396;
    wire N__29395;
    wire N__29394;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29371;
    wire N__29370;
    wire N__29369;
    wire N__29368;
    wire N__29367;
    wire N__29366;
    wire N__29365;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29357;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29316;
    wire N__29315;
    wire N__29312;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29291;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29209;
    wire N__29202;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29188;
    wire N__29185;
    wire N__29176;
    wire N__29173;
    wire N__29168;
    wire N__29165;
    wire N__29158;
    wire N__29155;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29137;
    wire N__29132;
    wire N__29127;
    wire N__29122;
    wire N__29117;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29053;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29014;
    wire N__29013;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29005;
    wire N__29004;
    wire N__29003;
    wire N__29002;
    wire N__29001;
    wire N__29000;
    wire N__28999;
    wire N__28998;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28978;
    wire N__28975;
    wire N__28974;
    wire N__28973;
    wire N__28970;
    wire N__28969;
    wire N__28968;
    wire N__28965;
    wire N__28960;
    wire N__28959;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28955;
    wire N__28954;
    wire N__28951;
    wire N__28950;
    wire N__28949;
    wire N__28946;
    wire N__28945;
    wire N__28944;
    wire N__28943;
    wire N__28942;
    wire N__28941;
    wire N__28940;
    wire N__28939;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28933;
    wire N__28932;
    wire N__28931;
    wire N__28930;
    wire N__28929;
    wire N__28928;
    wire N__28927;
    wire N__28926;
    wire N__28925;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28893;
    wire N__28890;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28870;
    wire N__28867;
    wire N__28858;
    wire N__28855;
    wire N__28850;
    wire N__28841;
    wire N__28828;
    wire N__28819;
    wire N__28814;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28781;
    wire N__28780;
    wire N__28779;
    wire N__28778;
    wire N__28775;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28767;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28749;
    wire N__28740;
    wire N__28733;
    wire N__28726;
    wire N__28723;
    wire N__28716;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28696;
    wire N__28691;
    wire N__28684;
    wire N__28677;
    wire N__28658;
    wire N__28657;
    wire N__28656;
    wire N__28655;
    wire N__28654;
    wire N__28653;
    wire N__28652;
    wire N__28651;
    wire N__28650;
    wire N__28649;
    wire N__28648;
    wire N__28647;
    wire N__28646;
    wire N__28645;
    wire N__28642;
    wire N__28641;
    wire N__28640;
    wire N__28639;
    wire N__28638;
    wire N__28637;
    wire N__28634;
    wire N__28633;
    wire N__28628;
    wire N__28623;
    wire N__28622;
    wire N__28621;
    wire N__28620;
    wire N__28619;
    wire N__28618;
    wire N__28617;
    wire N__28616;
    wire N__28615;
    wire N__28614;
    wire N__28613;
    wire N__28608;
    wire N__28603;
    wire N__28602;
    wire N__28601;
    wire N__28600;
    wire N__28599;
    wire N__28598;
    wire N__28593;
    wire N__28588;
    wire N__28587;
    wire N__28586;
    wire N__28585;
    wire N__28582;
    wire N__28577;
    wire N__28576;
    wire N__28575;
    wire N__28572;
    wire N__28563;
    wire N__28562;
    wire N__28561;
    wire N__28560;
    wire N__28559;
    wire N__28558;
    wire N__28557;
    wire N__28556;
    wire N__28551;
    wire N__28546;
    wire N__28545;
    wire N__28544;
    wire N__28539;
    wire N__28534;
    wire N__28529;
    wire N__28528;
    wire N__28527;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28511;
    wire N__28506;
    wire N__28503;
    wire N__28498;
    wire N__28495;
    wire N__28490;
    wire N__28485;
    wire N__28480;
    wire N__28475;
    wire N__28468;
    wire N__28461;
    wire N__28458;
    wire N__28453;
    wire N__28448;
    wire N__28443;
    wire N__28442;
    wire N__28441;
    wire N__28440;
    wire N__28437;
    wire N__28432;
    wire N__28429;
    wire N__28428;
    wire N__28427;
    wire N__28426;
    wire N__28425;
    wire N__28420;
    wire N__28415;
    wire N__28406;
    wire N__28401;
    wire N__28392;
    wire N__28385;
    wire N__28378;
    wire N__28373;
    wire N__28370;
    wire N__28365;
    wire N__28360;
    wire N__28353;
    wire N__28346;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28273;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28217;
    wire N__28216;
    wire N__28213;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28142;
    wire N__28141;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28112;
    wire N__28109;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28070;
    wire N__28069;
    wire N__28064;
    wire N__28061;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28037;
    wire N__28036;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28018;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27988;
    wire N__27985;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27950;
    wire N__27949;
    wire N__27944;
    wire N__27941;
    wire N__27940;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27869;
    wire N__27866;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27749;
    wire N__27748;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27716;
    wire N__27715;
    wire N__27710;
    wire N__27707;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27640;
    wire N__27637;
    wire N__27636;
    wire N__27633;
    wire N__27632;
    wire N__27631;
    wire N__27630;
    wire N__27629;
    wire N__27628;
    wire N__27625;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27611;
    wire N__27610;
    wire N__27609;
    wire N__27606;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27595;
    wire N__27594;
    wire N__27591;
    wire N__27590;
    wire N__27587;
    wire N__27582;
    wire N__27579;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27564;
    wire N__27559;
    wire N__27556;
    wire N__27551;
    wire N__27550;
    wire N__27545;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27513;
    wire N__27510;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27486;
    wire N__27479;
    wire N__27472;
    wire N__27461;
    wire N__27460;
    wire N__27457;
    wire N__27456;
    wire N__27455;
    wire N__27454;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27450;
    wire N__27449;
    wire N__27448;
    wire N__27447;
    wire N__27446;
    wire N__27445;
    wire N__27444;
    wire N__27443;
    wire N__27442;
    wire N__27441;
    wire N__27440;
    wire N__27439;
    wire N__27436;
    wire N__27435;
    wire N__27434;
    wire N__27433;
    wire N__27432;
    wire N__27431;
    wire N__27430;
    wire N__27429;
    wire N__27428;
    wire N__27425;
    wire N__27410;
    wire N__27395;
    wire N__27394;
    wire N__27393;
    wire N__27392;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27388;
    wire N__27387;
    wire N__27386;
    wire N__27385;
    wire N__27384;
    wire N__27381;
    wire N__27374;
    wire N__27371;
    wire N__27354;
    wire N__27347;
    wire N__27332;
    wire N__27327;
    wire N__27322;
    wire N__27321;
    wire N__27320;
    wire N__27317;
    wire N__27316;
    wire N__27315;
    wire N__27314;
    wire N__27313;
    wire N__27312;
    wire N__27309;
    wire N__27298;
    wire N__27295;
    wire N__27290;
    wire N__27289;
    wire N__27288;
    wire N__27287;
    wire N__27286;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27278;
    wire N__27277;
    wire N__27276;
    wire N__27275;
    wire N__27274;
    wire N__27273;
    wire N__27268;
    wire N__27263;
    wire N__27260;
    wire N__27253;
    wire N__27252;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27231;
    wire N__27226;
    wire N__27217;
    wire N__27212;
    wire N__27207;
    wire N__27206;
    wire N__27205;
    wire N__27200;
    wire N__27193;
    wire N__27192;
    wire N__27191;
    wire N__27188;
    wire N__27187;
    wire N__27186;
    wire N__27183;
    wire N__27178;
    wire N__27173;
    wire N__27170;
    wire N__27165;
    wire N__27160;
    wire N__27155;
    wire N__27152;
    wire N__27147;
    wire N__27142;
    wire N__27131;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26978;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26720;
    wire N__26717;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26624;
    wire N__26621;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26579;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26519;
    wire N__26516;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26447;
    wire N__26444;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26420;
    wire N__26419;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26233;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26189;
    wire N__26186;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26168;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26126;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26114;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26089;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26050;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25921;
    wire N__25918;
    wire N__25913;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25883;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25785;
    wire N__25784;
    wire N__25783;
    wire N__25782;
    wire N__25777;
    wire N__25774;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25763;
    wire N__25762;
    wire N__25761;
    wire N__25756;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25720;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25693;
    wire N__25690;
    wire N__25685;
    wire N__25680;
    wire N__25673;
    wire N__25670;
    wire N__25669;
    wire N__25668;
    wire N__25667;
    wire N__25662;
    wire N__25661;
    wire N__25660;
    wire N__25659;
    wire N__25658;
    wire N__25653;
    wire N__25650;
    wire N__25645;
    wire N__25640;
    wire N__25639;
    wire N__25638;
    wire N__25637;
    wire N__25636;
    wire N__25635;
    wire N__25632;
    wire N__25627;
    wire N__25624;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25609;
    wire N__25606;
    wire N__25605;
    wire N__25604;
    wire N__25603;
    wire N__25602;
    wire N__25601;
    wire N__25598;
    wire N__25593;
    wire N__25590;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25574;
    wire N__25571;
    wire N__25566;
    wire N__25561;
    wire N__25556;
    wire N__25541;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25504;
    wire N__25501;
    wire N__25498;
    wire N__25493;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25406;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25391;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25339;
    wire N__25336;
    wire N__25335;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25291;
    wire N__25288;
    wire N__25283;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25241;
    wire N__25238;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25220;
    wire N__25217;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25147;
    wire N__25144;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25129;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25034;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24952;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24917;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24866;
    wire N__24863;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24667;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24500;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24445;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24413;
    wire N__24410;
    wire N__24409;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24352;
    wire N__24349;
    wire N__24344;
    wire N__24341;
    wire N__24340;
    wire N__24339;
    wire N__24338;
    wire N__24337;
    wire N__24334;
    wire N__24333;
    wire N__24332;
    wire N__24331;
    wire N__24328;
    wire N__24327;
    wire N__24324;
    wire N__24323;
    wire N__24320;
    wire N__24319;
    wire N__24318;
    wire N__24317;
    wire N__24316;
    wire N__24315;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24309;
    wire N__24308;
    wire N__24301;
    wire N__24294;
    wire N__24293;
    wire N__24292;
    wire N__24291;
    wire N__24290;
    wire N__24289;
    wire N__24288;
    wire N__24279;
    wire N__24278;
    wire N__24277;
    wire N__24276;
    wire N__24275;
    wire N__24272;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24250;
    wire N__24245;
    wire N__24240;
    wire N__24237;
    wire N__24230;
    wire N__24227;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24203;
    wire N__24194;
    wire N__24187;
    wire N__24178;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24167;
    wire N__24166;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24162;
    wire N__24161;
    wire N__24156;
    wire N__24155;
    wire N__24154;
    wire N__24153;
    wire N__24148;
    wire N__24147;
    wire N__24144;
    wire N__24139;
    wire N__24136;
    wire N__24127;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24113;
    wire N__24112;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24098;
    wire N__24097;
    wire N__24096;
    wire N__24095;
    wire N__24094;
    wire N__24091;
    wire N__24086;
    wire N__24083;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24063;
    wire N__24054;
    wire N__24045;
    wire N__24036;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24014;
    wire N__24013;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23999;
    wire N__23994;
    wire N__23991;
    wire N__23990;
    wire N__23989;
    wire N__23988;
    wire N__23987;
    wire N__23986;
    wire N__23985;
    wire N__23982;
    wire N__23977;
    wire N__23976;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23927;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23908;
    wire N__23905;
    wire N__23894;
    wire N__23891;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23782;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23600;
    wire N__23597;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23534;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23486;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23462;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23411;
    wire N__23408;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23390;
    wire N__23387;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23375;
    wire N__23372;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23360;
    wire N__23359;
    wire N__23356;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23164;
    wire N__23163;
    wire N__23160;
    wire N__23159;
    wire N__23158;
    wire N__23155;
    wire N__23154;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23146;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23108;
    wire N__23107;
    wire N__23106;
    wire N__23105;
    wire N__23104;
    wire N__23103;
    wire N__23100;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23092;
    wire N__23089;
    wire N__23078;
    wire N__23071;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22979;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22949;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22913;
    wire N__22910;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22898;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22834;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22816;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22751;
    wire N__22748;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22652;
    wire N__22649;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22577;
    wire N__22576;
    wire N__22571;
    wire N__22568;
    wire N__22567;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22561;
    wire N__22560;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22524;
    wire N__22521;
    wire N__22516;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22502;
    wire N__22501;
    wire N__22498;
    wire N__22493;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22442;
    wire N__22439;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22388;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22376;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22294;
    wire N__22293;
    wire N__22292;
    wire N__22291;
    wire N__22290;
    wire N__22289;
    wire N__22288;
    wire N__22287;
    wire N__22286;
    wire N__22285;
    wire N__22284;
    wire N__22283;
    wire N__22280;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22272;
    wire N__22269;
    wire N__22268;
    wire N__22267;
    wire N__22266;
    wire N__22263;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22255;
    wire N__22252;
    wire N__22251;
    wire N__22248;
    wire N__22247;
    wire N__22246;
    wire N__22245;
    wire N__22242;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22234;
    wire N__22233;
    wire N__22232;
    wire N__22231;
    wire N__22230;
    wire N__22227;
    wire N__22210;
    wire N__22193;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22159;
    wire N__22156;
    wire N__22151;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22139;
    wire N__22138;
    wire N__22137;
    wire N__22136;
    wire N__22135;
    wire N__22134;
    wire N__22133;
    wire N__22132;
    wire N__22129;
    wire N__22124;
    wire N__22121;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22092;
    wire N__22089;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22071;
    wire N__22066;
    wire N__22063;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22045;
    wire N__22044;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22040;
    wire N__22039;
    wire N__22036;
    wire N__22031;
    wire N__22028;
    wire N__22019;
    wire N__22014;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21980;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21856;
    wire N__21855;
    wire N__21852;
    wire N__21847;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21836;
    wire N__21835;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21821;
    wire N__21818;
    wire N__21811;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21706;
    wire N__21703;
    wire N__21702;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21690;
    wire N__21687;
    wire N__21686;
    wire N__21685;
    wire N__21684;
    wire N__21683;
    wire N__21682;
    wire N__21677;
    wire N__21674;
    wire N__21669;
    wire N__21662;
    wire N__21655;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21580;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21548;
    wire N__21547;
    wire N__21546;
    wire N__21543;
    wire N__21538;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21517;
    wire N__21516;
    wire N__21509;
    wire N__21508;
    wire N__21507;
    wire N__21504;
    wire N__21499;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21457;
    wire N__21456;
    wire N__21455;
    wire N__21454;
    wire N__21453;
    wire N__21452;
    wire N__21449;
    wire N__21448;
    wire N__21447;
    wire N__21446;
    wire N__21445;
    wire N__21444;
    wire N__21443;
    wire N__21442;
    wire N__21441;
    wire N__21440;
    wire N__21439;
    wire N__21438;
    wire N__21437;
    wire N__21436;
    wire N__21433;
    wire N__21432;
    wire N__21429;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21411;
    wire N__21406;
    wire N__21403;
    wire N__21402;
    wire N__21401;
    wire N__21400;
    wire N__21399;
    wire N__21392;
    wire N__21391;
    wire N__21390;
    wire N__21389;
    wire N__21388;
    wire N__21383;
    wire N__21380;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21357;
    wire N__21356;
    wire N__21355;
    wire N__21350;
    wire N__21345;
    wire N__21342;
    wire N__21337;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21319;
    wire N__21316;
    wire N__21311;
    wire N__21306;
    wire N__21301;
    wire N__21296;
    wire N__21293;
    wire N__21284;
    wire N__21281;
    wire N__21274;
    wire N__21271;
    wire N__21260;
    wire N__21253;
    wire N__21250;
    wire N__21245;
    wire N__21244;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21226;
    wire N__21225;
    wire N__21224;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21216;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21212;
    wire N__21211;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21193;
    wire N__21190;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21182;
    wire N__21181;
    wire N__21180;
    wire N__21179;
    wire N__21176;
    wire N__21171;
    wire N__21164;
    wire N__21157;
    wire N__21152;
    wire N__21147;
    wire N__21144;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21107;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21083;
    wire N__21082;
    wire N__21081;
    wire N__21080;
    wire N__21079;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21061;
    wire N__21058;
    wire N__21047;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20998;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20980;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20965;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20857;
    wire N__20856;
    wire N__20855;
    wire N__20854;
    wire N__20853;
    wire N__20852;
    wire N__20851;
    wire N__20850;
    wire N__20849;
    wire N__20848;
    wire N__20847;
    wire N__20846;
    wire N__20843;
    wire N__20842;
    wire N__20841;
    wire N__20832;
    wire N__20831;
    wire N__20828;
    wire N__20813;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20794;
    wire N__20787;
    wire N__20782;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20735;
    wire N__20732;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20713;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20659;
    wire N__20658;
    wire N__20657;
    wire N__20648;
    wire N__20647;
    wire N__20646;
    wire N__20645;
    wire N__20644;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20640;
    wire N__20639;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20628;
    wire N__20627;
    wire N__20624;
    wire N__20609;
    wire N__20606;
    wire N__20597;
    wire N__20592;
    wire N__20587;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20542;
    wire N__20541;
    wire N__20540;
    wire N__20539;
    wire N__20536;
    wire N__20535;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20527;
    wire N__20524;
    wire N__20519;
    wire N__20514;
    wire N__20507;
    wire N__20502;
    wire N__20497;
    wire N__20494;
    wire N__20489;
    wire N__20486;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20467;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20440;
    wire N__20437;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20425;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20372;
    wire N__20369;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20332;
    wire N__20327;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20317;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20295;
    wire N__20288;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20189;
    wire N__20186;
    wire N__20185;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20056;
    wire N__20053;
    wire N__20052;
    wire N__20051;
    wire N__20050;
    wire N__20047;
    wire N__20046;
    wire N__20045;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20014;
    wire N__20011;
    wire N__20004;
    wire N__20001;
    wire N__19996;
    wire N__19993;
    wire N__19988;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19963;
    wire N__19960;
    wire N__19959;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19951;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19947;
    wire N__19946;
    wire N__19945;
    wire N__19944;
    wire N__19943;
    wire N__19940;
    wire N__19939;
    wire N__19938;
    wire N__19937;
    wire N__19936;
    wire N__19933;
    wire N__19932;
    wire N__19931;
    wire N__19926;
    wire N__19919;
    wire N__19918;
    wire N__19917;
    wire N__19914;
    wire N__19909;
    wire N__19904;
    wire N__19903;
    wire N__19902;
    wire N__19901;
    wire N__19898;
    wire N__19887;
    wire N__19880;
    wire N__19875;
    wire N__19872;
    wire N__19871;
    wire N__19870;
    wire N__19869;
    wire N__19866;
    wire N__19859;
    wire N__19852;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19819;
    wire N__19816;
    wire N__19809;
    wire N__19806;
    wire N__19799;
    wire N__19798;
    wire N__19797;
    wire N__19796;
    wire N__19795;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19784;
    wire N__19783;
    wire N__19782;
    wire N__19781;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19777;
    wire N__19776;
    wire N__19771;
    wire N__19768;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19751;
    wire N__19744;
    wire N__19743;
    wire N__19740;
    wire N__19739;
    wire N__19734;
    wire N__19729;
    wire N__19722;
    wire N__19717;
    wire N__19714;
    wire N__19709;
    wire N__19706;
    wire N__19701;
    wire N__19698;
    wire N__19691;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19651;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19632;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19618;
    wire N__19617;
    wire N__19614;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19586;
    wire N__19581;
    wire N__19580;
    wire N__19579;
    wire N__19578;
    wire N__19577;
    wire N__19572;
    wire N__19569;
    wire N__19564;
    wire N__19563;
    wire N__19558;
    wire N__19557;
    wire N__19556;
    wire N__19555;
    wire N__19552;
    wire N__19551;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19515;
    wire N__19508;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19486;
    wire N__19483;
    wire N__19482;
    wire N__19479;
    wire N__19478;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19472;
    wire N__19471;
    wire N__19468;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19444;
    wire N__19441;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19420;
    wire N__19415;
    wire N__19412;
    wire N__19407;
    wire N__19404;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19375;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19330;
    wire N__19325;
    wire N__19322;
    wire N__19321;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19283;
    wire N__19280;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19258;
    wire N__19255;
    wire N__19250;
    wire N__19247;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19236;
    wire N__19235;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19221;
    wire N__19218;
    wire N__19213;
    wire N__19208;
    wire N__19207;
    wire N__19206;
    wire N__19205;
    wire N__19204;
    wire N__19203;
    wire N__19202;
    wire N__19201;
    wire N__19200;
    wire N__19195;
    wire N__19190;
    wire N__19189;
    wire N__19188;
    wire N__19187;
    wire N__19186;
    wire N__19181;
    wire N__19180;
    wire N__19177;
    wire N__19172;
    wire N__19167;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19153;
    wire N__19152;
    wire N__19147;
    wire N__19144;
    wire N__19137;
    wire N__19134;
    wire N__19129;
    wire N__19126;
    wire N__19121;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19069;
    wire N__19068;
    wire N__19067;
    wire N__19066;
    wire N__19065;
    wire N__19062;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19058;
    wire N__19057;
    wire N__19056;
    wire N__19053;
    wire N__19046;
    wire N__19043;
    wire N__19042;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19018;
    wire N__19013;
    wire N__19010;
    wire N__19009;
    wire N__19006;
    wire N__19005;
    wire N__19002;
    wire N__19001;
    wire N__19000;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18980;
    wire N__18977;
    wire N__18972;
    wire N__18969;
    wire N__18964;
    wire N__18961;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18935;
    wire N__18932;
    wire N__18931;
    wire N__18930;
    wire N__18929;
    wire N__18928;
    wire N__18927;
    wire N__18926;
    wire N__18925;
    wire N__18922;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18914;
    wire N__18913;
    wire N__18912;
    wire N__18909;
    wire N__18908;
    wire N__18903;
    wire N__18898;
    wire N__18895;
    wire N__18890;
    wire N__18885;
    wire N__18884;
    wire N__18883;
    wire N__18880;
    wire N__18875;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18863;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18841;
    wire N__18836;
    wire N__18833;
    wire N__18828;
    wire N__18821;
    wire N__18812;
    wire N__18811;
    wire N__18806;
    wire N__18803;
    wire N__18802;
    wire N__18801;
    wire N__18798;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18784;
    wire N__18783;
    wire N__18778;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18766;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18750;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18724;
    wire N__18719;
    wire N__18716;
    wire N__18715;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18571;
    wire N__18568;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18461;
    wire N__18458;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18446;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18418;
    wire N__18413;
    wire N__18410;
    wire N__18409;
    wire N__18406;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18371;
    wire N__18370;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18349;
    wire N__18344;
    wire N__18341;
    wire N__18340;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18307;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18244;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18199;
    wire N__18194;
    wire N__18193;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18172;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18160;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18122;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18076;
    wire N__18073;
    wire N__18070;
    wire N__18067;
    wire N__18064;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18043;
    wire N__18042;
    wire N__18039;
    wire N__18034;
    wire N__18033;
    wire N__18030;
    wire N__18029;
    wire N__18026;
    wire N__18025;
    wire N__18024;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18004;
    wire N__17993;
    wire N__17992;
    wire N__17991;
    wire N__17990;
    wire N__17989;
    wire N__17988;
    wire N__17985;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17974;
    wire N__17971;
    wire N__17964;
    wire N__17961;
    wire N__17960;
    wire N__17959;
    wire N__17954;
    wire N__17951;
    wire N__17946;
    wire N__17943;
    wire N__17938;
    wire N__17931;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17890;
    wire N__17887;
    wire N__17886;
    wire N__17883;
    wire N__17882;
    wire N__17881;
    wire N__17872;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17861;
    wire N__17860;
    wire N__17859;
    wire N__17858;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17850;
    wire N__17849;
    wire N__17846;
    wire N__17841;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17815;
    wire N__17804;
    wire N__17803;
    wire N__17802;
    wire N__17801;
    wire N__17800;
    wire N__17799;
    wire N__17798;
    wire N__17795;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17776;
    wire N__17775;
    wire N__17774;
    wire N__17773;
    wire N__17772;
    wire N__17771;
    wire N__17768;
    wire N__17763;
    wire N__17760;
    wire N__17755;
    wire N__17746;
    wire N__17739;
    wire N__17732;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17640;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17609;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17585;
    wire N__17582;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17531;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17443;
    wire N__17442;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17430;
    wire N__17429;
    wire N__17426;
    wire N__17425;
    wire N__17420;
    wire N__17417;
    wire N__17416;
    wire N__17415;
    wire N__17414;
    wire N__17413;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17405;
    wire N__17404;
    wire N__17403;
    wire N__17402;
    wire N__17401;
    wire N__17400;
    wire N__17395;
    wire N__17394;
    wire N__17391;
    wire N__17390;
    wire N__17387;
    wire N__17380;
    wire N__17379;
    wire N__17374;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17341;
    wire N__17340;
    wire N__17339;
    wire N__17336;
    wire N__17331;
    wire N__17322;
    wire N__17315;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17285;
    wire N__17282;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17260;
    wire N__17259;
    wire N__17256;
    wire N__17255;
    wire N__17252;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17234;
    wire N__17231;
    wire N__17230;
    wire N__17227;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17211;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17156;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17142;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17128;
    wire N__17127;
    wire N__17126;
    wire N__17125;
    wire N__17124;
    wire N__17123;
    wire N__17122;
    wire N__17121;
    wire N__17110;
    wire N__17103;
    wire N__17102;
    wire N__17101;
    wire N__17100;
    wire N__17097;
    wire N__17092;
    wire N__17089;
    wire N__17084;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17003;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16989;
    wire N__16984;
    wire N__16981;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16861;
    wire N__16858;
    wire N__16855;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16824;
    wire N__16823;
    wire N__16822;
    wire N__16821;
    wire N__16816;
    wire N__16811;
    wire N__16806;
    wire N__16799;
    wire N__16798;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16757;
    wire N__16756;
    wire N__16753;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16694;
    wire N__16691;
    wire N__16686;
    wire N__16685;
    wire N__16684;
    wire N__16683;
    wire N__16680;
    wire N__16679;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16648;
    wire N__16645;
    wire N__16634;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16623;
    wire N__16620;
    wire N__16619;
    wire N__16616;
    wire N__16615;
    wire N__16610;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16594;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16578;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16552;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16510;
    wire N__16507;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16495;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16483;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16468;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16441;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16393;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16361;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16295;
    wire N__16292;
    wire N__16291;
    wire N__16290;
    wire N__16289;
    wire N__16288;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16280;
    wire N__16279;
    wire N__16278;
    wire N__16277;
    wire N__16276;
    wire N__16275;
    wire N__16272;
    wire N__16271;
    wire N__16270;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16246;
    wire N__16237;
    wire N__16234;
    wire N__16233;
    wire N__16232;
    wire N__16231;
    wire N__16230;
    wire N__16229;
    wire N__16228;
    wire N__16227;
    wire N__16226;
    wire N__16225;
    wire N__16224;
    wire N__16223;
    wire N__16222;
    wire N__16221;
    wire N__16220;
    wire N__16219;
    wire N__16218;
    wire N__16217;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16112;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16012;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15976;
    wire N__15971;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15959;
    wire N__15958;
    wire N__15957;
    wire N__15956;
    wire N__15955;
    wire N__15954;
    wire N__15949;
    wire N__15946;
    wire N__15941;
    wire N__15940;
    wire N__15939;
    wire N__15938;
    wire N__15937;
    wire N__15936;
    wire N__15935;
    wire N__15934;
    wire N__15933;
    wire N__15932;
    wire N__15929;
    wire N__15928;
    wire N__15927;
    wire N__15926;
    wire N__15921;
    wire N__15918;
    wire N__15913;
    wire N__15910;
    wire N__15903;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15869;
    wire N__15866;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15826;
    wire N__15823;
    wire N__15820;
    wire N__15817;
    wire N__15814;
    wire N__15811;
    wire N__15808;
    wire N__15803;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15763;
    wire N__15762;
    wire N__15759;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15729;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15611;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15450;
    wire N__15449;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15441;
    wire N__15438;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15403;
    wire N__15400;
    wire N__15393;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15370;
    wire N__15369;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15350;
    wire N__15349;
    wire N__15348;
    wire N__15347;
    wire N__15342;
    wire N__15337;
    wire N__15332;
    wire N__15331;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15176;
    wire N__15167;
    wire N__15166;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15158;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15144;
    wire N__15141;
    wire N__15136;
    wire N__15133;
    wire N__15128;
    wire N__15125;
    wire N__15122;
    wire N__15113;
    wire N__15110;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15102;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15049;
    wire N__15046;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15035;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15020;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14974;
    wire N__14973;
    wire N__14970;
    wire N__14969;
    wire N__14968;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14932;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14824;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14809;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14791;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14662;
    wire N__14661;
    wire N__14660;
    wire N__14659;
    wire N__14658;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14611;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14578;
    wire N__14577;
    wire N__14574;
    wire N__14573;
    wire N__14570;
    wire N__14569;
    wire N__14568;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14560;
    wire N__14559;
    wire N__14556;
    wire N__14555;
    wire N__14554;
    wire N__14553;
    wire N__14548;
    wire N__14541;
    wire N__14538;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14516;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14491;
    wire N__14488;
    wire N__14487;
    wire N__14486;
    wire N__14485;
    wire N__14484;
    wire N__14481;
    wire N__14478;
    wire N__14473;
    wire N__14468;
    wire N__14465;
    wire N__14456;
    wire N__14455;
    wire N__14454;
    wire N__14449;
    wire N__14446;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14366;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14354;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14330;
    wire N__14327;
    wire N__14326;
    wire N__14325;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14294;
    wire N__14293;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14275;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14240;
    wire N__14237;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14225;
    wire N__14222;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14124;
    wire N__14123;
    wire N__14122;
    wire N__14121;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14075;
    wire N__14074;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14059;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13941;
    wire N__13940;
    wire N__13939;
    wire N__13938;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13879;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13831;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13730;
    wire N__13729;
    wire N__13728;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13682;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13657;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13636;
    wire N__13633;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13597;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13586;
    wire N__13585;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13561;
    wire N__13558;
    wire N__13555;
    wire N__13552;
    wire N__13549;
    wire N__13546;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13501;
    wire N__13500;
    wire N__13497;
    wire N__13492;
    wire N__13487;
    wire N__13486;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13459;
    wire N__13456;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13429;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13405;
    wire N__13402;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13366;
    wire N__13363;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13355;
    wire N__13352;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13338;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13324;
    wire N__13319;
    wire N__13316;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13304;
    wire N__13301;
    wire N__13300;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13279;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13261;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13222;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13210;
    wire N__13205;
    wire N__13202;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13037;
    wire N__13036;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13006;
    wire N__13003;
    wire N__13000;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12979;
    wire N__12976;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12944;
    wire N__12943;
    wire N__12940;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12898;
    wire N__12895;
    wire N__12890;
    wire N__12885;
    wire N__12878;
    wire N__12875;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12790;
    wire N__12787;
    wire N__12784;
    wire N__12781;
    wire N__12778;
    wire N__12775;
    wire N__12772;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12757;
    wire N__12754;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12733;
    wire N__12730;
    wire N__12727;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12692;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12645;
    wire N__12640;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12536;
    wire N__12533;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12499;
    wire N__12498;
    wire N__12495;
    wire N__12490;
    wire N__12487;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12382;
    wire N__12379;
    wire N__12376;
    wire N__12371;
    wire N__12368;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12355;
    wire N__12350;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12332;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12283;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12264;
    wire N__12263;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12249;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12177;
    wire N__12176;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12162;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12103;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12040;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12028;
    wire N__12023;
    wire VCCG0;
    wire GNDG0;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_5 ;
    wire \processor_zipi8.flags_i.un5_shift_carry_value_cascade_ ;
    wire \processor_zipi8.flags_i.shift_carry_value_1_0_0_cascade_ ;
    wire \processor_zipi8.stack_i.data_out_ram_0 ;
    wire \processor_zipi8.shadow_carry_flag ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI88F42_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV3DI8_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIM5NP1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINR4G8_7 ;
    wire \processor_zipi8.port_id_7_cascade_ ;
    wire \processor_zipi8.port_id_7 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_7 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_7 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_7_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_7 ;
    wire \processor_zipi8.stack_memory_5 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_5 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_5_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_5 ;
    wire \processor_zipi8.port_id_5_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_5 ;
    wire \processor_zipi8.port_id_5 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_5 ;
    wire \processor_zipi8.stack_memory_9 ;
    wire \processor_zipi8.stack_memory_4 ;
    wire \processor_zipi8.stack_memory_8 ;
    wire \processor_zipi8.stack_memory_10 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_9 ;
    wire \processor_zipi8.sy_5 ;
    wire \processor_zipi8.sy_7 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_8 ;
    wire \processor_zipi8.pc_vector_8_cascade_ ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_9_cascade_ ;
    wire address_9;
    wire \processor_zipi8.program_counter_i.un380_half_pc_cascade_ ;
    wire \processor_zipi8.program_counter_i.half_pc_0_10_cascade_ ;
    wire address_10;
    wire \processor_zipi8.return_vector_10 ;
    wire \processor_zipi8.program_counter_i.un395_half_pcZ0 ;
    wire \processor_zipi8.program_counter_i.carry_pc_46_7 ;
    wire \processor_zipi8.pc_vector_8 ;
    wire \processor_zipi8.program_counter_i.carry_pc_46_7_cascade_ ;
    wire address_8;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_8 ;
    wire \processor_zipi8.flags_i.zero_flag_3_cascade_ ;
    wire \processor_zipi8.shadow_zero_flag ;
    wire \processor_zipi8.alu_result_7 ;
    wire \processor_zipi8.alu_result_6_cascade_ ;
    wire \processor_zipi8.flags_i.zero_flag_3_0_5 ;
    wire \processor_zipi8.alu_result_5 ;
    wire \processor_zipi8.stack_i.stack_zero_flag ;
    wire \processor_zipi8.stack_i.shadow_zero_value ;
    wire \processor_zipi8.alu_result_3 ;
    wire \processor_zipi8.flags_i.m82_1_cascade_ ;
    wire \processor_zipi8.flags_i.m82_1 ;
    wire \processor_zipi8.zero_flag_RNIJSPM4 ;
    wire \processor_zipi8.flags_i.N_55 ;
    wire \processor_zipi8.flags_i.m61_ns_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIK2TR1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_7 ;
    wire \processor_zipi8.spm_data_5 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_6 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_6_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_6 ;
    wire \processor_zipi8.sy_6 ;
    wire \processor_zipi8.port_id_6_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_6 ;
    wire \processor_zipi8.port_id_6 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_6 ;
    wire \processor_zipi8.stack_memory_6 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_6 ;
    wire \processor_zipi8.flags_i.N_125_mux_cascade_ ;
    wire \processor_zipi8.stack_i.stack_bit ;
    wire \processor_zipi8.run ;
    wire BTN1_c;
    wire \processor_zipi8.stack_memory_2 ;
    wire \processor_zipi8.special_bit ;
    wire \processor_zipi8.state_machine_i.bram_enable ;
    wire \processor_zipi8.stack_memory_11 ;
    wire \processor_zipi8.flags_i.N_37 ;
    wire \processor_zipi8.stack_memory_7 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_7 ;
    wire \processor_zipi8.stack_memory_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_155 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_195_cascade_ ;
    wire address_6;
    wire address_4;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_4 ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_4_cascade_ ;
    wire \processor_zipi8.program_counter_i.carry_pc_28_4_cascade_ ;
    wire \processor_zipi8.program_counter_i.carry_pc_34_5 ;
    wire \processor_zipi8.pc_vector_6 ;
    wire \processor_zipi8.program_counter_i.carry_pc_34_5_cascade_ ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_6 ;
    wire \processor_zipi8.program_counter_i.carry_pc_40_6 ;
    wire \processor_zipi8.pc_vector_7 ;
    wire \processor_zipi8.program_counter_i.carry_pc_40_6_cascade_ ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_7 ;
    wire address_7;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_5 ;
    wire \processor_zipi8.pc_vector_5 ;
    wire \processor_zipi8.program_counter_i.carry_pc_28_4 ;
    wire address_5;
    wire \processor_zipi8.return_vector_11 ;
    wire \processor_zipi8.program_counter_i.un3_half_pcZ0_cascade_ ;
    wire \processor_zipi8.program_counter_i.half_pc_0_10 ;
    wire \processor_zipi8.program_counter_i.un431_half_pc ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_11_cascade_ ;
    wire \processor_zipi8.address_11 ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_9 ;
    wire \processor_zipi8.pc_vector_9 ;
    wire \processor_zipi8.program_counter_i.carry_pc_52_8 ;
    wire \processor_zipi8.program_counter_i.carry_pc_58_9 ;
    wire \processor_zipi8.flags_i.m49_ns_1 ;
    wire \processor_zipi8.flags_i.N_50_cascade_ ;
    wire \processor_zipi8.flags_i.N_51_cascade_ ;
    wire \processor_zipi8.flags_i.N_123_mux ;
    wire \processor_zipi8.flags_i.N_45 ;
    wire \processor_zipi8.flags_i.m91_amZ0_cascade_ ;
    wire \processor_zipi8.flags_i.m25_ns_1_cascade_ ;
    wire \processor_zipi8.flags_i.N_26_0_cascade_ ;
    wire \processor_zipi8.flags_i.N_27_0 ;
    wire \processor_zipi8.flags_i.m20_ns_1_cascade_ ;
    wire \processor_zipi8.flags_i.N_21_0 ;
    wire \processor_zipi8.flags_i.N_1235_cascade_ ;
    wire \processor_zipi8.flags_i.zero_flag_RNI89VZ0Z91 ;
    wire \processor_zipi8.flags_i.N_1239 ;
    wire \processor_zipi8.flags_i.N_124_mux ;
    wire \processor_zipi8.flags_i.N_1241_cascade_ ;
    wire \processor_zipi8.zero_flag_RNIDS654 ;
    wire \processor_zipi8.stack_pointer_1 ;
    wire \processor_zipi8.flags_i.m75_amZ0 ;
    wire \processor_zipi8.flags_i.m75_amZ0_cascade_ ;
    wire \processor_zipi8.flags_i.zero_flag_RNI3VCZ0Z94 ;
    wire \processor_zipi8.zero_flag_RNI5GK75 ;
    wire \processor_zipi8.flags_i.N_1241 ;
    wire \processor_zipi8.stack_pointer_0 ;
    wire \processor_zipi8.stack_pointer_2 ;
    wire \processor_zipi8.flags_i.N_54 ;
    wire \processor_zipi8.flags_i.m68_ns_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_6 ;
    wire \processor_zipi8.spm_data_6 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe8 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe11 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212_cascade_ ;
    wire \processor_zipi8.shift_rotate_result_6 ;
    wire \processor_zipi8.shift_rotate_result_5 ;
    wire \processor_zipi8.port_id_2_cascade_ ;
    wire \processor_zipi8.port_id_2 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_2 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_2 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_2_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_2 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_2 ;
    wire \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_0_cascade_ ;
    wire instruction_2;
    wire \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_1_cascade_ ;
    wire \processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_0 ;
    wire address_2;
    wire \processor_zipi8.stack_pointer_4 ;
    wire \processor_zipi8.flags_i.N_34 ;
    wire \processor_zipi8.port_id_0_cascade_ ;
    wire \processor_zipi8.stack_memory_0 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_0 ;
    wire \processor_zipi8.pc_vector_0 ;
    wire \processor_zipi8.pc_vector_0_cascade_ ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_0 ;
    wire \processor_zipi8.flags_i.i14_mux ;
    wire \processor_zipi8.flags_i.i14_mux_0 ;
    wire \processor_zipi8.zero_flag_RNIC4FP9 ;
    wire \processor_zipi8.program_counter_i.t_state_0_1 ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_1_cascade_ ;
    wire \processor_zipi8.program_counter_i.half_pc_0_1_cascade_ ;
    wire address_1;
    wire \processor_zipi8.program_counter_i.half_pc_0_0 ;
    wire address_0;
    wire \processor_zipi8.zero_flag_RNIL8RB5 ;
    wire \processor_zipi8.program_counter_i.half_pc_0_1 ;
    wire \processor_zipi8.program_counter_i.carry_pc_4_0 ;
    wire \processor_zipi8.program_counter_i.carry_pc_22_3 ;
    wire \processor_zipi8.pc_vector_2 ;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_2 ;
    wire \processor_zipi8.program_counter_i.half_pc_0_2 ;
    wire \processor_zipi8.program_counter_i.un3_half_pcZ0 ;
    wire \processor_zipi8.program_counter_i.half_pc_0_3 ;
    wire \processor_zipi8.un16_alu_mux_sel_value_cascade_ ;
    wire \processor_zipi8.decode4_strobes_enables_i.un23_flag_enable_type ;
    wire \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_1_cascade_ ;
    wire \processor_zipi8.shift_rotate_result_2 ;
    wire \processor_zipi8.spm_data_2 ;
    wire \processor_zipi8.register_bank_control_i.un31_regbank_type_3_cascade_ ;
    wire \processor_zipi8.register_bank_control_i.un31_regbank_type ;
    wire \processor_zipi8.shift_rotate_result_0 ;
    wire \processor_zipi8.spm_data_0 ;
    wire \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_0_cascade_ ;
    wire \processor_zipi8.pc_mode_2_0_0 ;
    wire \processor_zipi8.decode4_pc_statck_i.un3_pc_modeZ0 ;
    wire \processor_zipi8.N_17_0 ;
    wire bram_enable_g;
    wire \processor_zipi8.flags_i.m104Z0Z_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI44F42_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIK4HN1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNII1NP1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIGUSR1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7B4G8_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe13 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe15 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe9 ;
    wire \processor_zipi8.sx_7 ;
    wire \processor_zipi8.sx_6 ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6 ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_7 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_6 ;
    wire \processor_zipi8.flags_i.carry_flag_value_1_1_cascade_ ;
    wire \processor_zipi8.flags_i.parity_4 ;
    wire \processor_zipi8.flags_i.carry_flag_RNOZ0Z_1 ;
    wire \processor_zipi8.flags_i.arith_carryZ0 ;
    wire \processor_zipi8.flags_i.shift_carryZ0 ;
    wire \processor_zipi8.flags_i.carry_flag_value_1_0_0 ;
    wire \processor_zipi8.decode4_pc_statck_i.N_22_0 ;
    wire \processor_zipi8.register_bank_control_i.un17_regbank_type_1 ;
    wire \processor_zipi8.flags_i.un17_carry_flag_value_0 ;
    wire \processor_zipi8.alu_mux_sel_value_1 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2 ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_0_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_0_cascade_ ;
    wire \processor_zipi8.port_id_0 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_0 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4Z0Z_0 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0 ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1 ;
    wire instruction_0;
    wire \processor_zipi8.register_bank_control_i.un1_bank_value ;
    wire \processor_zipi8.register_bank_control_i.bank_0_1_cascade_ ;
    wire \processor_zipi8.sy_4 ;
    wire \processor_zipi8.stack_i.stack_bank ;
    wire \processor_zipi8.shadow_bank ;
    wire \processor_zipi8.un16_alu_mux_sel_value ;
    wire \processor_zipi8.un4_arith_logical_sel_cascade_ ;
    wire \processor_zipi8.flags_i.carry_flag_value_1_0 ;
    wire \processor_zipi8.internal_reset ;
    wire \processor_zipi8.flags_i.N_69 ;
    wire \processor_zipi8.stack_pointer_3 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_3_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_3 ;
    wire \processor_zipi8.port_id_3_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_3 ;
    wire \processor_zipi8.port_id_3 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_3 ;
    wire instruction_3;
    wire \processor_zipi8.pc_vector_3 ;
    wire \processor_zipi8.pc_mode_2 ;
    wire \processor_zipi8.pc_mode_1 ;
    wire address_3;
    wire \processor_zipi8.program_counter_i.half_pc_0_0_3 ;
    wire \processor_zipi8.arith_carry_in_0 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0 ;
    wire \processor_zipi8.returni_type_o_2 ;
    wire \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_3 ;
    wire \processor_zipi8.decode4_strobes_enables_i.un9_flag_enable_type_cascade_ ;
    wire \processor_zipi8.decode4_strobes_enables_i.flag_enable_type_0_cascade_ ;
    wire \processor_zipi8.flag_enable ;
    wire \processor_zipi8.decode4_strobes_enables_i.spm_enable_value_1 ;
    wire \processor_zipi8.spm_enable ;
    wire \processor_zipi8.flags_i.use_zero_flagZ0 ;
    wire \processor_zipi8.alu_result_0_cascade_ ;
    wire \processor_zipi8.zero_flag ;
    wire \processor_zipi8.carry_flag ;
    wire \processor_zipi8.N_11_0 ;
    wire \processor_zipi8.alu_result_1 ;
    wire \processor_zipi8.alu_result_2_cascade_ ;
    wire \processor_zipi8.flags_i.zero_flag_3_0_0 ;
    wire \processor_zipi8.flags_i.zero_flag_3_0_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe12 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_bm_1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_179 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_am_1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_4_cascade_ ;
    wire \processor_zipi8.shift_rotate_result_4 ;
    wire \processor_zipi8.spm_data_4 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4 ;
    wire \processor_zipi8.shift_rotate_result_1 ;
    wire \processor_zipi8.spm_data_1 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3 ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2 ;
    wire \processor_zipi8.decode4_strobes_enables_i.un8_register_enable_type ;
    wire \processor_zipi8.t_state_1 ;
    wire \processor_zipi8.decode4_strobes_enables_i.register_enable_type_0_cascade_ ;
    wire instruction_17;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_22_3 ;
    wire \processor_zipi8.sx_5 ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_34_5 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_5 ;
    wire \processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4 ;
    wire \processor_zipi8.flags_i.parity_5 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_1_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tzZ0Z_4 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_4_cascade_ ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_4 ;
    wire \processor_zipi8.port_id_4 ;
    wire \processor_zipi8.arith_logical_sel_1 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_4 ;
    wire \processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical ;
    wire \processor_zipi8.un4_arith_logical_sel ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1Z0Z_1 ;
    wire \processor_zipi8.arith_and_logic_operations_i.N_773_tz ;
    wire \processor_zipi8.arith_logical_sel_1_0_0 ;
    wire \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_4 ;
    wire instruction_14;
    wire \processor_zipi8.arith_logical_sel_1_0_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_3 ;
    wire \processor_zipi8.sy_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_bm_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI8OGN1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_am_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIONE42_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI6LMP1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI4ISR1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINP2G8_3_cascade_ ;
    wire \processor_zipi8.sx_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6 ;
    wire \processor_zipi8.alu_result_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI43VU1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIGMK32_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIO8HN1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNICBE42_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIQ8MP1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIO5SR1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI781G8_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209 ;
    wire \processor_zipi8.register_enable ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNISBGN1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram15_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram8_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram9_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram11_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram10_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram12_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram13_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_7 ;
    wire \processor_zipi8.port_id_1 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_1 ;
    wire instruction_1;
    wire \processor_zipi8.pc_vector_1 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_4 ;
    wire instruction_12;
    wire \processor_zipi8.pc_vector_4 ;
    wire instruction_13;
    wire \processor_zipi8.sx_0 ;
    wire LED1_c;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_119_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_95 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_151 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_175 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_191_cascade_ ;
    wire \processor_zipi8.sx_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNII4IQ1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI4AK32_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIOMUU1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI8MSR1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIAPMP1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFIBI8_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7A3G8_4_cascade_ ;
    wire \processor_zipi8.sx_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNISRE42_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI4KGN1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIKJE42_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI0ESR1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI2HMP1_2 ;
    wire \processor_zipi8.sx_addr_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI792G8_2_cascade_ ;
    wire \processor_zipi8.sx_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_0 ;
    wire \processor_zipi8.shift_rotate_result_3 ;
    wire \processor_zipi8.spm_data_3 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_7 ;
    wire CONSTANT_ONE_NET;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNICIK32_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFJCI8_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI0VUU1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIQCIQ1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_243_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_299 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_315 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_219 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_275 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIUGIQ1_7 ;
    wire \processor_zipi8.shift_rotate_result_7 ;
    wire \processor_zipi8.spm_data_7 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNICSGN1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1211 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_0 ;
    wire \processor_zipi8.sy_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_1 ;
    wire \processor_zipi8.sy_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe23 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_123 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_99_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_5 ;
    wire \processor_zipi8.stack_memory_3 ;
    wire \processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_3 ;
    wire instruction_16;
    wire instruction_15;
    wire \processor_zipi8.un28_carry_flag_value_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_6_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNISIMM1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe28 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI86UU1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNI2KHQ1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFG9I8_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_0_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIKPJ32_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI4QLM1_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe16 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_5_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram7_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_2_cascade_ ;
    wire instruction_7;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_2_cascade_ ;
    wire \processor_zipi8.bank ;
    wire \processor_zipi8.sy_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe29 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe27 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_4_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIKAMM1_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_271 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_311 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram30_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_295 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_1_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_215 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_239 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIASHQ1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIC2MM1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFHAI8_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIS1K32_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIGEUU1_2_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI06K32_3_cascade_ ;
    wire instruction_10;
    wire instruction_11;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIE0IQ1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV1BI8_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIG6MM1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram19_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIKIUU1_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram17_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_3_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram31_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe24 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe25 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_5 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_6 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe26 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_7_cascade_ ;
    wire instruction_5;
    wire instruction_6;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram25_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram24_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_7_cascade_ ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI0NMM1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram26_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram27_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_7 ;
    wire instruction_9;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram28_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram29_7 ;
    wire instruction_8;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_3 ;
    wire \processor_zipi8.arith_logical_result_5 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5 ;
    wire \processor_zipi8.arith_logical_result_6 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_6 ;
    wire \processor_zipi8.arith_logical_result_7 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram20_4 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20 ;
    wire \processor_zipi8.arith_logical_result_0 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0 ;
    wire \processor_zipi8.arith_logical_result_1 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_1 ;
    wire \processor_zipi8.arith_logical_result_2 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_2 ;
    wire \processor_zipi8.arith_logical_result_3 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram23_3 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3 ;
    wire instruction_4;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_3 ;
    wire \processor_zipi8.alu_mux_sel_1 ;
    wire \processor_zipi8.arith_logical_result_4 ;
    wire \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ;
    wire \processor_zipi8.alu_mux_sel_0 ;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.ram22_4 ;
    wire CLK_3P3_MHZ_c_g;
    wire \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22 ;
    wire _gnd_net_;

    defparam \test_program.Ram2048x2_inst3_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst3_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_F=256'b0010011000100001000000100010000000000010000000000000011000100100001001100000000000000000001000000000000000000001000000000000000000100000001000000010000000100000000000010000100100001000000010000000100000001000000111000001100100011000001010000001100000011001;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_E=256'b0000110000001100000010000000100000001001000000000001010000010100000000010000000100000101000001000000000000000000000001000000010000000100000001000000000100000100001001010000010100000100000001000000010100000000000000000000000000100110001001100000001100000011;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_D=256'b0000011000000110001000110010000100000000001000000010001000100000000000100000101100101000000010110001111000011111001010110000100100001000000010000010101100101001000010110000100100001010001010000010101000100000001000100010000100000000000000010010000100100001;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_C=256'b0010001000100010000000010000000100100001001000010000000000000000001000000010000000000000001000000010000000000000001000000001000000000000000100010010100100111000000010000001100000101000001110000000100000011001000010000011100100101000001010010001100100011001;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_B=256'b0001000000010000000100010000000100010001000100000000001000000010001000000010000000000000000000010001000000000001000000010000000000001000000010000001000100011000000010010000100000001000000010000000000000001000000000000000000000000000000000000000000000000000;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_A=256'b0000000000000001000110000001000000010000000000010001000000010001000100000000000100010010000110110000000000000001000010000000000000001000000010010001100000001001000010000000100100001000000010000001100000011001000010000000100100000000000000010000000000000000;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_9=256'b0000000100000000000000000000000000000000000000000000000000000001000100000001000000010010000000000001100100010000000100100000100000011000000010010001000000001000000000100000000100000100001000000001001000110000000101110011000000010010001000000000101000100000;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_8=256'b0001001000110001000000100011000100100010001000000010100000100000001000000000000000100010000000100010000000000000001010010000000000001000001010000000100000101000000011010010110000001000001010000000110000101100000010010010100000000000001000000000000000100001;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_7=256'b0000010000100000000100000010000000000100001000010000000000100000000000000010000000010000001000010000100000100000000000000010100000001010001110100000100000101000000000000010100100000000001001010000010000100101000011000010010100100100001001000010110000100101;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_6=256'b0010010000000101001011000000010100110100000001010010010000011001000100000011010000010100001001000001010000110100000001000010010000000100001001000000010000110000000101100010001000000100001100010000010000100001000101000011100100001100001010010000100000101001;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_5=256'b0000100000111000000110000010110100001100001111010000110000101000000100000011000100000010001000010000000000100101000001000011000100010000001000010000001000110111000001100010001100010100000101100000000000011010000001100000100100001000000111010001010000001101;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_4=256'b0000010000010101000000000000000100010100000100010000000100010100000001010000000100000001000100000001001100000101000001000001000000000011000000000001001100010001000001000011010000000001000000100000000100110011000100000010001000000001001100100000000100100010;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_3=256'b0000001000110001000100000011000000010010001100100000000100100000000000010010001000000000001000000000000100100011000010100011000000000001001100000000000000100000000100000000001000010001000100010000000000000000000000010000001100000000000000010001000000000001;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_2=256'b0000000000000001000000000000000100000000000000010000000000001001000000000000000100000010000000110000100000000011000000000000000100010010000000110000000000000001000010000000000101010000000000010101001000000011011100000101000100000100000000010000000000000001;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_1=256'b0000001001000011010000000000000100010000010000010001000000010001010000100100011100000000000000010000000000000001000000000100000101000010001000110000000001100001000000000010000101000000011000000000001000100010000000000010000000000000011000000100000000100000;
    defparam \test_program.Ram2048x2_inst3_physical .INIT_0=256'b0000001001100010000010000010000001000000011000000000000100100001000000100010001000000000011000000100000000000000000000010100000100000000000000000100010001000000000000000100000000000001000000000000010001000100010001000000111000000100010001000000010000000100;
    SB_RAM40_4K \test_program.Ram2048x2_inst3_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,instruction_7,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,instruction_6,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__12595,N__12757,N__13003,N__14194,N__13798,N__14011,N__13648,N__17698,N__15292,N__15682,N__15505}),
            .WADDR({N__12592,N__12754,N__13000,N__14185,N__13795,N__14002,N__13645,N__17695,N__15277,N__15679,N__15508}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45}),
            .RCLKE(N__16223),
            .RCLK(N__33659),
            .RE(N__22529),
            .WCLKE(N__16222),
            .WCLK(N__33658),
            .WE());
    defparam \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical .WRITE_MODE=0;
    defparam \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \processor_zipi8.spm_with_output_reg_i.spm_ram.ram_s_ram_s_0_0_physical  (
            .RDATA({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,\processor_zipi8.spm_data_7 ,\processor_zipi8.spm_data_6 ,\processor_zipi8.spm_data_5 ,\processor_zipi8.spm_data_4 ,\processor_zipi8.spm_data_3 ,\processor_zipi8.spm_data_2 ,\processor_zipi8.spm_data_1 ,\processor_zipi8.spm_data_0 }),
            .RADDR({dangling_wire_54,dangling_wire_55,dangling_wire_56,N__12197,N__13366,N__12284,N__19246,N__17186,N__15049,N__21569,N__16840}),
            .WADDR({dangling_wire_57,dangling_wire_58,dangling_wire_59,N__12196,N__13370,N__12283,N__19247,N__17185,N__15050,N__21565,N__16841}),
            .MASK({dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75}),
            .WDATA({dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,N__16701,N__16632,N__18803,N__21860,N__20056,N__22049,N__21707,N__21112}),
            .RCLKE(),
            .RCLK(N__33619),
            .RE(N__22562),
            .WCLKE(N__17477),
            .WCLK(N__33618),
            .WE(N__22560));
    defparam \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical .WRITE_MODE=0;
    defparam \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \processor_zipi8.stack_i.stack_ram.ram_s_ram_s_0_0_physical  (
            .RDATA({\processor_zipi8.stack_memory_11 ,\processor_zipi8.stack_memory_10 ,\processor_zipi8.stack_memory_9 ,\processor_zipi8.stack_memory_8 ,\processor_zipi8.stack_memory_7 ,\processor_zipi8.stack_memory_6 ,\processor_zipi8.stack_memory_5 ,\processor_zipi8.stack_memory_4 ,\processor_zipi8.stack_memory_3 ,\processor_zipi8.stack_memory_2 ,\processor_zipi8.stack_memory_1 ,\processor_zipi8.stack_memory_0 ,\processor_zipi8.stack_i.stack_bit ,\processor_zipi8.stack_i.stack_bank ,\processor_zipi8.stack_i.stack_zero_flag ,\processor_zipi8.stack_i.data_out_ram_0 }),
            .RADDR({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,N__15779,N__15386,N__14603,N__13076,N__14690}),
            .WADDR({dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,N__15166,N__17261,N__14501,N__14675,N__14582}),
            .MASK({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111}),
            .WDATA({N__14402,N__12543,N__12692,N__12944,N__14124,N__13740,N__13941,N__13596,N__17608,N__15204,N__15630,N__15450,N__13502,N__25637,N__18047,N__17992}),
            .RCLKE(),
            .RCLK(N__33617),
            .RE(N__22563),
            .WCLKE(N__19070),
            .WCLK(N__33620),
            .WE(N__22561));
    defparam \test_program.Ram2048x2_inst6_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst6_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_F=256'b0000101000011100000011100001100100001000001111010010110000011001000010000001110100111111000111110001101000111100001111100001110100011110001111010001010000011101000111100001111100011110000111110001111000011111000010110000101100011000000111110001101000101110;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_E=256'b0001111000111011001110100011111100100010001001110011011000111011001010110010111000101110001010100010101000101111001011110010101100101110001010110000101100101110001011100010101000101110000010110011101000111110001010000011111100011110001110010000101100101110;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_D=256'b0000111000101001001010000000101100001010001011110010000000001111000011100010110000101010000010100001101000101001001011010001111000111110001111110010111100001100001011110010110000001100001011010010011100000111001001100000111000001110001011110010011100001110;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_C=256'b0010110000001111000001010010111000101111000011100000011000101111001011100000111000000110001011100010111000001110001101100001111000011110001111100011111100010110000111100011111100111110000111110001111000111110001111100001111000101110000111110000111100101110;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_B=256'b0011010000101111001011110010111000001111001011100011110000111111000111010011111100111110000111100000111000001111001111110011111000111110001101110010111100101110001101110011111000011110000111110001111000011110000111100001111000011110000111100001011000011110;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_A=256'b0001101000011110000101100000111100001110001111100011011000001111000011100010111000000100001011110011110000111110001111100011011100111110001111100010101000101111001111100011111000111110001111110010111000101110000111100001111100010110000111100001111000011111;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_9=256'b0001111100011110000111110001111100011010000111110001111000011110001111100010111100101100001011010010111000100110001111000010110100100110001111100011110000101111001111100011110000111000001110110011111000101101001000010011101000101111001011010010101000100001;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_8=256'b0010100000101001001000100010101100101010000110110011101100010011001110110001101100110000000110110010100000011011001111110001011000111110000111110010101000101011001010110010101000101010001010110010101000101011001010100010101100100110001011110010101100101110;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_7=256'b0010111100101011001111100010111100111010001111110011111000111111001111100011111100101101001011100011111000110111001111100011111100110100001011110010110000111111001010100010111100101110001011110010111000101111001011100010011100101110000011110010011000001111;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_6=256'b0010111000001111001011100000011100101110000011110011011000001011000010100001111100100110001000110010011000100011001001100010001100100110001100110011011000100011001001000010001100110100001000110010001000110011001010100010001100101010001010110010111000111111;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_5=256'b0011101000101111001011100010101100111010001010110010101000111011001001000010111100101010001011110010111000111001001110100010111100101110001011110011110000101011001010100001100100001010001010010000110000000111000010110001110000010101000010100000100000001001;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_4=256'b0001100100001000000011000001110100000001000011000000110000001000000010000001110000011100000011000000111000001000000110000000111100001110000111000000111000001100001011000000111100001010001110000011110000101110001011100010110100111100001011100010111000111100;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_3=256'b0011011000100101001011000011111100101110001011000010010000101110001011100010000000100101001011100010101000100100001001100010110000111000001111100010111100111010001110100010110100110000001100100010001000110011001100100011000100110011001100010011000100100011;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_2=256'b0011001101110001011000010001001100010011011100110001111100111011000111010001110100001001000111010001000100011001000110010001001100010001000010010000101100010011000100010001101100111001000010110000000100111001001110110000101100011001001110110011100101111111;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_1=256'b0111100100101101001011110011101101111101001011110010100101101111001111010011100100111111001110110001100101111011010011010011111100111001001111010111111100111011001000010110011100101101001011110010110100101101001000110110111101101101001000110010000100101111;
    defparam \test_program.Ram2048x2_inst6_physical .INIT_0=256'b0110110100100101001001110110111100101100001111110011110000101110001011000111110101110110001001110010010000110111011101000010011000100100011101110010000000110011001101000011001100110110011101000111010100110010000111010011101001011101001110100001110101111010;
    SB_RAM40_4K \test_program.Ram2048x2_inst6_physical  (
            .RDATA({dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,instruction_13,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,instruction_12,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .RADDR({N__12559,N__12721,N__12967,N__14158,N__13762,N__13975,N__13612,N__17662,N__15256,N__15646,N__15469}),
            .WADDR({N__12556,N__12718,N__12964,N__14149,N__13759,N__13966,N__13609,N__17659,N__15241,N__15643,N__15472}),
            .MASK({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141}),
            .WDATA({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157}),
            .RCLKE(N__16225),
            .RCLK(N__33694),
            .RE(N__22556),
            .WCLKE(N__16224),
            .WCLK(N__33693),
            .WE());
    defparam \test_program.Ram2048x2_inst1_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst1_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_F=256'b0010000000101000000000000000100100000000001000000010010000000110000000100000001000000001001000010000000000100010000000000010001000100000001000000010000000110000000010000011101000001000001110100000101000111000000010110010100100001000000010000000100000001010;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_E=256'b0000100000001010000100000000001000000000001010100000000000100000000000000010000100000100001001000000000000000000000011100000111000001110000010100000101000001010000010110000101100001011000101000000001000000000001000100000000000110100001101000000000000000011;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_D=256'b0000000000000000000000010000010100000010000000000010000000100000000010110000101000101010001111100000111000011011001111010010100000111110000110000000110100001000001011000000100100100001001000000010100100001101000000010010010000001010000001010000000000010100;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_C=256'b0000101000100010000000000000000000001001001000110000000100000010000011010000011100000101000001110010110100010101001001010011010100001100000101000010110000110100000011110000111000101110000010100000111100001010000011100010101000001110000010010000111000001100;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_B=256'b0010111000001100001111100001110000011111000110010001111100001010001111010010100100001101000000100000100000000011000110010010011000011000001011100010100100001100001000000000010100000001000000000001100100011001000110110001001100011011000100110001001100010011;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_A=256'b0001101000000010000001100010010000001111000001000010011100000000000111110001000000010111000100100010110100110000001010010001111000101001000011100010100100001010001010010001101000001000001110000000100100101000001111010001110000111101000011000011110100001110;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_9=256'b0011110100001110001111000000101000101000000110100010100100110000001010000010000000111000000100000011000000010000001110000001110000100001000001000001100100111100000110010010011000011011001000010001110000100110000100000011000000011100000101000000000000011000;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_8=256'b0001100000000000000100000001000000001000000000000000001000001000000110000001000000000010000000100000100000000100000011000000111000011000000110100001100000101110000110010010101000011001001011000001100000001000000110000000110100011100000011000001000100001011;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_7=256'b0001000000111010000101000011111000000000001010100001000100010000000000000000000000000011000000000000000000000001001110000011100000110010001100100010000100000000001010000000101100100100000001110010010100000111000001010010111100001100000001000000010000000101;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_6=256'b0000110000000101000001000001110000001000000000110001000000000011000110010001001000101000001000100011100000111000001010000000000000111000000010000011100000000000001010100000101100001001001100010011100000101000001110000011111000101100000011100011110100001110;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_5=256'b0011100000001010001010010000100100001100001011010001110000101100000111000011110100000001001010010001010100001101000100000000100000000111000010010001001000000011000100000010010100010001000100100000010100000101000110100000100000010001000000010000110000001100;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_4=256'b0000000000000000000101000000010000010001000100010000100000001000000110010000000100011000000000010000101000000111000110000000000000010110000010010001111000111111000010010010100000001000000110110011110000101101001011100010010000101100000100010010010100011010;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_3=256'b0011011000000010001111000001100000011011001101100000000100110101000011000011110000000001001100000000100100011011000001110000011000011011000100010000010100001010001100000011101000111111000100010011111100011001001011010000001100111101000110010001110100110001;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_2=256'b0001111100111000000011010100000000011111000111000000111100001100001010000000001100100010000000010011011000010011001011000000000100110100000100100010110000000000001101000111001000111100001100000000010100000011011001010110010100010001001001110111100100101000;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_1=256'b0110110100001010001010010000100000111001010110100110010000001001010100000111111100000000001010010100000000001011010000000000000000110000001100100010110000100010011100000000000001111101010010010011000100000010011100010000001001010001001001010001000100100000;
    defparam \test_program.Ram2048x2_inst1_physical .INIT_0=256'b0101010100100011010100000011001001001100010001000001110000010100010011010000001001011001000101100000100000001100000111000001000001101100001010000110100001100010001110000011110001111001001100000111100000001001000110000000100101010000000000110101100000000001;
    SB_RAM40_4K \test_program.Ram2048x2_inst1_physical  (
            .RDATA({dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,instruction_3,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,instruction_2,dangling_wire_169,dangling_wire_170,dangling_wire_171}),
            .RADDR({N__12619,N__12781,N__13027,N__14218,N__13822,N__14035,N__13672,N__17722,N__15314,N__15706,N__15529}),
            .WADDR({N__12616,N__12778,N__13024,N__14209,N__13819,N__14026,N__13669,N__17719,N__15301,N__15703,N__15532}),
            .MASK({dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187}),
            .WDATA({dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203}),
            .RCLKE(N__16231),
            .RCLK(N__33696),
            .RE(N__22501),
            .WCLKE(N__16230),
            .WCLK(N__33695),
            .WE());
    defparam \test_program.Ram2048x2_inst4_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst4_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_F=256'b0011101000000011000111100001110100101000000010110000111000010000001001110000110000000101000101000000101000101001001111110001010000010100001010110010000100010101000010110000100000011110000101100001010100001000000000010001011000011001000110010011100000010001;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_E=256'b0001010100001010000100100011000100001011000000100000010000000000000000000001011000000110000010000000101000010010000011010000100000000100000100110000001100001001000011100011001000001100001010010010100000011011000010100010000000100100001010100000001000000100;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_D=256'b0011110000111010000110000010001000100010000111000000001000100011001110000001101000011110001001110010010100001011000001100010000000001011001011110000110000100010000100100011110000110111000000010000110100110101000000000010011000110100000100010001010000100110;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_C=256'b0000001000100011001100000001010000010100001000000010010000010111000000100010000100010010001100110001010000100001000101000010011100110011000101010000111000101011001001000001110000011000001000100001101000111100000001100010001100000101001011010000100000110110;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_B=256'b0010111100001001000001100011110000001010000000100001101100111111000101010000000100010100001111000001100000000011001110100001100000111010001011110000110000011000000011000010011000001010000100010011101000101111001111000001000100001100001011110000001000010001;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_A=256'b0011001100100011001000000000000000010000000001100000011000100001001001100001011000100010001000110001000000010100000111000010100100110100000111100011101000100001000110100001101000010000001001010010010000011010000011100000010100001010001110100011000000001101;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_9=256'b0011110000110010000011110000110100000011001100100011000000001100000011000000011000001110001110010010101100001101001010100010101000011110000001100000110000101001001110000000011000001000000111010000010000100010001101000001011000100101001101110001101100011100;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_8=256'b0001001100100001001100010001010000100000000000100000100000101100000000000001001000100010001101100010000000000001000010000010110000000000000100100000001100001001000011100011001000111001000010000011010100110010000000110000100100001010001100100011000000000000;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_7=256'b0011010100111010000010100000000100001011001010100010010000010101001001000011101100001010000001000000101100101000000011110001111000001110001000110010100000010101001110000011100100011100000001110000111000111001001010100000111100110000000100010001010000100111;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_6=256'b0000011000010001001010100010111100100000000100010000010000100011000101100000010100110110001001110001010000001001000000000010011100110010000010010010011000100111000101100000101100000000001001010000000000011011000111000010100100100100000000010011000000101001;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_5=256'b0000100000000001000111000010100100100100000001010010010000111001000110000000000100000000001000110011010000001011001010100010000100011000000010110000011000100011000001000011101100111100000001110000101000101001000110000000101000101110001000000011110000001111;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_4=256'b0000110000100100000010000001101100110000001000000010010000000010000100000010100000001000000000100011110000101010001000100000000100000000001110100001000000000010000000100010100100111000000000100000111000001000000100000010011100100100000010100010110000110110;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_3=256'b0000100100000010000010110011010100111100000000110010011000100100000011000000101000000000001001100010100000001010001001000010001100010110000100100001111000100010000010010000101100011010001100100011101100001110001111000010001100011100000111100000101000100000;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_2=256'b0010100000001110010011000010001000101110011111000110110001001010010010100001011000000010011000000010001000010010011010000110110001000100000000000000111001101110001010000000101000001010011011000101010000010000010101100011011000110100001010100101101000010100;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_1=256'b0000100000101000011101100001001000100000001011100000001001000000010001000011100000101010000001100110100000011010001001100010010001000100000110000000111000100010001010000100001001101010001100000001100000000100010100100011001000101100000010100110001000110000;
    defparam \test_program.Ram2048x2_inst4_physical .INIT_0=256'b0001100000001000000100100111001001110000000101100010111000100100010111000001110000001110001000110100110100001110000010100010000000111000010111000110110000100011000011010000101001001000001100100011111000001100011111100011100000001000000001100000000001110010;
    SB_RAM40_4K \test_program.Ram2048x2_inst4_physical  (
            .RDATA({dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,instruction_9,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,instruction_8,dangling_wire_215,dangling_wire_216,dangling_wire_217}),
            .RADDR({N__12583,N__12745,N__12991,N__14182,N__13786,N__13999,N__13636,N__17686,N__15280,N__15670,N__15493}),
            .WADDR({N__12580,N__12742,N__12988,N__14173,N__13783,N__13990,N__13633,N__17683,N__15265,N__15667,N__15496}),
            .MASK({dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .WDATA({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .RCLKE(N__16218),
            .RCLK(N__33657),
            .RE(N__22530),
            .WCLKE(N__16219),
            .WCLK(N__33660),
            .WE());
    defparam \test_program.Ram2048x2_inst7_physical .INIT_0=256'b0010010100111001011011110111110100101100001001000010110000101100001011000010100000100110001010000011010000011000001001000000100001110100010110100010001000011010001101000001110000110000000111100011011000011100000101000001010000011110000101100101110001011100;
    defparam \test_program.Ram2048x2_inst7_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst7_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_F=256'b0000101000001011000010110000101100000010000000100000000000000101000001010001010100010100000100100011000000110111000100110001000100110011001100110001001100010011000100100011100100010010001110010001001100111001000000100011100000000001000010100000001000011011;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_E=256'b0001001100101011001100110010101100100010001100110010001000101011001011110011111000101011001111110010111000111110001010100011100000101010001110000000111100011101000010100001100000001010001111000010011000000100001000000000011100000000000000010000000000110000;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_D=256'b0000010000010010000000110011011100100011001100000000000000110110001000000011110000000000001110000010000000101010000101100001111000100110001011000000010000011010001001010001100000000101000111010000010000010100000001000011110000101110001111000000011000011100;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_C=256'b0000110000110100001001000011111000001111001111100010011100111111000011100001011100100110001111110000111000011011000101100010101100111110001001100001011100100110001111100010110000011110000011010011111000101100000111100000110000001110000111000010111000101000;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_B=256'b0010110000001010001011100000000000001111001000000011110100010001001111000001001000011110000000100001111000000010001111100000001000110110000010100010111000001010001111110000101000010111001000110001011000100011000111100010000100011110001000010001001000101101;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_A=256'b0001101000101100000001100011100100011110001100000000011000001000000011100000100000000100000010000011110000110010001101100011101000111110001010100011101000101110001111100010101000111110001010100010111000101010000111100010101000011110001010100001111000100000;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_9=256'b0001111000100000000111100010000000011010001001000001111000100100001011100000010000101101000001110010011000001101001011000001111100111110000111000010010000010100001111000000010000111000001001000010110000101001001100100011111100101001001000100010000100100100;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_8=256'b0010100000101100001000000010110000001000000101010001001100010100000110110001110000000000000011010000100100000110000101100000001000011110000010100010101100011010001010100001101100101011000110110010101100011010001010100001101000101110000111110010101000010001;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_7=256'b0010101100010000001011110000010000111010000100000011101000010000001110110000000100111000000000110011001100001001001110110010100000101000001110000011000000100010001000100011001000101010001101100010101000110110001000100011011000001010000111100000001000011110;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_6=256'b0000101000010110000000100001011000001010000011000000001000001000000111100001010000100010000010000010001000001000001000100000100000100010000010000010001000001000001000000000100000100000000010100011001000111010001000100010101000101010001010100010111000101110;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_5=256'b0010101000101010001010100010101000101010001010100011101000111010001011000010110000101000001000000010100000100000001011100010010000101110001000000010100000100000000110000011000000101000000000100000011000101110000010000010101000001010001010110000000100100011;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_4=256'b0000100000100010000111010011011100000000001010100000100000101010000011000010111000001100001010100000100000101010000011100010111000011100001110000000110000100110000010100000001000101000001001100010111000000010001011000000010000101110000001100011110000011100;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_3=256'b0010010000001110001101100001011000101100000001100010011000010110001000000001010000100110000100100010010000011000001011000000110000101010000000100010101000001001001011010010110100110010001111100011001000111100001100000010110000110001001011110010001100101111;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_2=256'b0011000101111101000000110100111101010011000111010001001101010001000011010110000100001101011010010001000101100101000100010110011100000001011101010001001101111101000110010110110100001001001001010011000100111101000010110000110100111001001010010011100100001001;
    defparam \test_program.Ram2048x2_inst7_physical .INIT_1=256'b0010100100001001001111110001100100101101000011010110110101010101001110010001000100111111000100010000110100000001000010010000000100111001001000010011101100101101011001010111110100100101001100010010100100110001001000110011000100100001001101010010010100110101;
    SB_RAM40_4K \test_program.Ram2048x2_inst7_physical  (
            .RDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,instruction_15,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,instruction_14,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RADDR({N__12547,N__12709,N__12955,N__14146,N__13750,N__13963,N__13600,N__17650,N__15244,N__15634,N__15457}),
            .WADDR({N__12544,N__12706,N__12952,N__14137,N__13747,N__13954,N__13597,N__17647,N__15228,N__15631,N__15460}),
            .MASK({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279}),
            .WDATA({dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295}),
            .RCLKE(N__16229),
            .RCLK(N__33707),
            .RE(N__22567),
            .WCLKE(N__16228),
            .WCLK(N__33706),
            .WE());
    defparam \test_program.Ram2048x2_inst2_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst2_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_F=256'b0000101000100011000010100010000000000000000000100010011000000100000000000010001000000001000100010000000000010001001000000001000000100010001100100000101000110000000010100001100000001010000110000000100000011010000110010001101100101000000010000001100000001011;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_E=256'b0001110000001110000010000011001000001000001000100001010000110110000010010010001000001100001000110000110000100010000001000010100000000100001010000000000000001000000001010000110000100100000010000010000000000000000000000010000000100010001001000000001000000010;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_D=256'b0000011000000000001000010000000100000000000000000000100000000000001010010000101100101111001010110001110000101111001011000010110100001101000011010010110000001101000011000000110100101100001000100000000000101000000000010010000100001000001010010010000000000001;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_C=256'b0000101100101011000000000010000100001000001010100010100000000010000011000010101000000000000000100000110000001010001000000010101000001000001010110000000000000011001010000000100000001000000010000010100100001001001010010010100100001000000010010001100000101000;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_B=256'b0010000100100001001100000010000000010001000100010000001000010010001000000011000000100001001000110011010000000011001000010001001100100001000100110001100100111011000110010010101100011000000010100000100000011010000000000001000000000000000100000000000000010000;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_A=256'b0000100000011001000001000000000000001101000010010000010000100000000111010000100100010110000100110011110100001001001111000000001100101101000010110011100000001010001111010000101100111101000010110011110100011011000110000000111100010001000001110001000000000101;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_9=256'b0001000000000101000100000000010000010000000000000001000100000101001000000000010000110000000001000011100100011100001010100001110000101001000011010011100000001100001100010001011100010100000100000001110000011010000100000001000100011000000110000001000000001000;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_8=256'b0001100000011011000010010000000000001000001010000001000000011000001110010010100100100010000010100000100000101000000101000001001000111100001011100000100000101010000011000010101000001000001010100000110000101010000010010010101000000100001000100000000100100001;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_7=256'b0000000000000000000001000000000000010000000100000001000000000001000000000000000000010001000000010001000000011000000110000000100000011010000010100000100100001000000011010000101000000101000001100000010100000110000001000000111000001101001011100000010100000110;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_6=256'b0010110100101111001001010000111000011101001010000001000000010000001110010011100000000101000101000000010100010000000000010001010000000001000000000001010100000100000001110001001100010000000001000000000000100011000011000011001100011000001011100000110000101010;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_5=256'b0001100100101010000011010011101000011101001010110000100100101110000001010011000000010001001100000000001100100100000100110010000000000001001100100000011100110010000001100000001100000010000101000000110000001000000010100000100000011110000010000000110100011001;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_4=256'b0000000000010100000001000000000100000000000100000000100000010100000010010000000100011100000000010000101000010110000010000000001100001010000001010000011000010010001101000000001000000100000000110001010000100000000001000011000000000100001000010000111000100001;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_3=256'b0001011000100011000101000011001000000100001100000000011000100000000011010010100000000011001010010000101100101011000101100011001000011100001110000000111100100101001011100000001000110001000100000010000000000010001100110001001100110010000000110010000000000011;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_2=256'b0011001000010011011000000000001100010010000000110001111000011111000000100000000100001010000000110001000000000001000110000001000100000010000000110000100000000011000100000001001101100000000000010000001001000010001110000100001000111100001100100011000000011000;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_1=256'b0111011000011110001001000101101001100000000010100011010000010100001100100100001000110100010101100000010000000010010000000000000000010010011000100101000000111110000000000010001000000101011001010100001100100011000000010010001101000001001011100000000101101001;
    defparam \test_program.Ram2048x2_inst2_physical .INIT_0=256'b0000011101101110000001010010011000001100011010100100010101101000000100100010111001000100001000100011010001000010001000010101010000010000001001000000010001100100000100000010000000010000001000000101010000100100000111000100100000010000000001000001000000001000;
    SB_RAM40_4K \test_program.Ram2048x2_inst2_physical  (
            .RDATA({dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,instruction_5,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,instruction_4,dangling_wire_307,dangling_wire_308,dangling_wire_309}),
            .RADDR({N__12607,N__12769,N__13015,N__14206,N__13810,N__14023,N__13660,N__17710,N__15304,N__15694,N__15517}),
            .WADDR({N__12604,N__12766,N__13012,N__14197,N__13807,N__14014,N__13657,N__17707,N__15289,N__15691,N__15520}),
            .MASK({dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325}),
            .WDATA({dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341}),
            .RCLKE(N__16227),
            .RCLK(N__33676),
            .RE(N__22502),
            .WCLKE(N__16226),
            .WCLK(N__33675),
            .WE());
    defparam \test_program.Ram2048x2_inst8_physical .INIT_0=256'b0110101101011000001001010101000001100100000000000011110100000000001010100100000001110000000110000000000001001000010100010101100000000010010010000101011000001000000101000000110000010111010011100101000100001110000100010100010001010011010001000001100101000100;
    defparam \test_program.Ram2048x2_inst8_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst8_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_F=256'b0010100000000010000011010000001000000000001010100010011100001100000100110010100000110010001010100001011000101010001100110010111000010001000011100011000100001110000100000010010000010001001001000001000100100100000000000010010000000010000000000000001000000000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_E=256'b0010011100000000001000110000000000101010000000000010111100000100001010110001000100101110000101010010101000010001001011000001000100101100000101010000100100010000000011010001000000001100000101010000000000011000000001010001100000000111000010000010000100011100;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_D=256'b0000011100011111001000000011110000000000000110010010010000111001000001110001010000100100001100000001011000010011001001010000000000100100000000010000000100010000000000010001000100000100000100010010110000010000001011010011000000001100000100010010010100010000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_C=256'b0010010000110001000011110001000000101111001100010000011000010001001001100011000100001110000100010010101000010001001000100010000100000110000000000010111000101000000001000000000000100101001000000000010100000000001001000000000000110100001000010001000100000000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_B=256'b0001000000000001000100010000000000110001000000010001000000100001000100100010000000000011001100000000001000110001000000110000000000001010000010010001001100001000000000110000100100000010001000010000001000100001000000000010000100000000001000010000110000100101;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_A=256'b0000110000100000000100010011000000100001000000000011100000000000000110010000000000010000001000000011001100000000001110100000100000100011000100000010011000010000001000110000000000100010000000000011001100000000000000100010000000000011001000000000000000100000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_9=256'b0000000100100000000000000010000100000100001000010000010100100000000101010000000100010100000000010001110100001000000101010001000000000101000000000001010000010000000001110000000000100000000000000011101100010010001000010001000100110000000000010011100000000101;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_8=256'b0011100000000100001100000000010000010001001001000001100100100100000110010010010000000001001101000000001000110100000010110010100000000011001000010000011000010001000001110001000100000110000100000000011000010000000001100001000000000111000100000000000100010001;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_7=256'b0000010000010001000101000000000100010000000000000001000000000100000000010001010000000001000101010000100000001100001000000000110000110001000111000010001100010100001000110001010000100011000100000010001100010000001010110001000000001011001100000000001100110000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_6=256'b0000001100110000000010110011000000001001001000000001010100110100000000010010000000000001000111000001000100001100000000010000110000000001000111000001000100001100000000010001110000010011000111000010001100011100001111110000100000100111000000000010011100010000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_5=256'b0011001100000000001001110001000000110111000100000010011100010000001101010000000000100001000000000010010100010100001100010000000000100001000100000011010100010000001001110011000000010111001000100000110100101000000000110011001000010101001000010000010000110011;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_4=256'b0001010100110011000001000011001100011001001000110000110100100110000010010011001000011001001000100000111100110110000110000011000000001011001100000001011100100010001000000010000000000011001100100001000100000000000001100001001000010101000100000000111100010000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_3=256'b0001011000010010000001000000000000010111000000100000010100010000000011110001011000000001000101000000101100011100000001110000001000000001000000000000110100000101001110100001001000100001000011000010000000001100001000100000110000100011000011100011000100001100;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_2=256'b0111001100001110011000010100110000010001011011000001010101100100000000110111010000001011011101000000001101100100000010110110010000010011011101000000100101101100000000010110010000110001001101000000101101000100011010010010010000001101001000000000100101000000;
    defparam \test_program.Ram2048x2_inst8_physical .INIT_1=256'b0101101100010000000011010100010001011001010001000000000101000100010101110000010000010001000001000000000101010100010000010001010000100011010001000110110101000100001000010101000001100001000100000010001100010100001000010101010001101101000101000010000101010000;
    SB_RAM40_4K \test_program.Ram2048x2_inst8_physical  (
            .RDATA({dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,instruction_17,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,dangling_wire_352,instruction_16,dangling_wire_353,dangling_wire_354,dangling_wire_355}),
            .RADDR({N__12536,N__12691,N__12939,N__14122,N__13729,N__13939,N__13585,N__17639,N__15234,N__15610,N__15448}),
            .WADDR({N__12532,N__12699,N__12951,N__14121,N__13728,N__13938,N__13584,N__17620,N__15214,N__15609,N__15437}),
            .MASK({dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371}),
            .WDATA({dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387}),
            .RCLKE(N__16217),
            .RCLK(N__33629),
            .RE(N__22568),
            .WCLKE(N__16216),
            .WCLK(N__33628),
            .WE());
    defparam \test_program.Ram2048x2_inst5_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst5_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_F=256'b0001100000001001001110000000100100111000000110010001100000111000001010000000110100001000001011010011100000000001000010000011010100101000000101010000100000010101001010000001110100101000000010000010100000001001001010000000100100111100000100010011100000010001;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_E=256'b0001100000010001000111000001000100010000000000010000000000000010000000000000001000000001000000100000000100000010000000000000000100000000000010010000000000001001000000000000100000000001000010100000000100001010000000000000101000110000001010000001010000001010;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_D=256'b0010000000110000000001110011000000000101000100100000000100010010000000000000100000000000000010110000000000011001000100100000110000110000001001110011001000100100001000100011010000100010001101010000001000110101000001100011000000000110000000010000011000100000;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_C=256'b0001011000100111000001000001010000000100001101000000010000010101000001000011000100000000000000010000000000000111000000000000011100000000000000110000000000010011000010010001000000001000001101000000100000010100000110000000110100001000001011110000110000011010;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_B=256'b0000110000011011000011000001001000001100000101100001111000010111000111000001110100011100000111000001110000011001000110000001100000010000000100010000000000011010000000000000101000100000000011110000000000101111000000000010110100000000001111010000000000110001;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_A=256'b0000000000010001000001000001001000000100000000100000010000110011001001000011001000100110001101110001010000010100000101000001010100011100000101000001100000010001000110000011000000011000001110110000100000111010000010000000101100001000000011100000100000000101;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_9=256'b0000100000000100000010010011010000001001001110000000110000111010000010000001111000001000000111110000000100010110000000000001111000000000001010100000001000111001000000000010100000000110000010010000010000010000000100100001010000000010000101010000011000100001;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_8=256'b0000011000100001000001100010000100000110001000000001011000100000000101100010000000010110000000100001010000000001000101000000000000010100000000000000000000000101000000000000000000000000000001110000000000001011000000000011111100000100001110100000010000110000;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_7=256'b0000000000110001001001000001000100110100000000010011000000001111001100000000111100110000001011100011000000100111000100000000101100000010000110110001000000001001000000000001100100000000001111010000000000111101000000000011010100000000001001110000000000100011;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_6=256'b0000000000100011000000000000001100010000000000010000000000010001000100000000010100011000001001010010100000000111001110000000011100111000000001110010100000010011001110100010001100101000001100010001100000000001000000000000000100010000000000010001000000000001;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_5=256'b0000000000110001000100000010000100000000001110010001000000101001001000000000100100110000000000010011000000000001001000000001000100110000001000010010001000111011000100000010100100100000001010010011000000100001001100000010100000100000000110000011001000001001;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_4=256'b0010001000011000001100100000100100000010001000000001001000100000000100100010000000000010001100000001000000000000000000010001100000010000000010000000010000000000000101010010000000110100001000000000000000010000000101010000100000000100000110000001010000001000;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_3=256'b0000010100111100000101010010110000000100001011000001010000100101001100000000000000110000000000000011000000000000001100000000000000100000001100010011000000101000000001000001100100010100000010000001010000001001000101000000100100010100001010000000010000111100;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_2=256'b0001010000101100000101000110110001110100001011000011000001101000000100000100100000010000010000000001010001000000000101000000000000000100001100000001010000100010000101000010111001000100001111100101010000010100000101000011011001110000001100100101000000010010;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_1=256'b0000000001010000010000000001101000000000010110100100000000100010000100000010000001010000001000100111000000100010001100000110101001010000000010000001000001001010010000000000111000000000000011100100000000101000010000000010001000000000011100100100000000110110;
    defparam \test_program.Ram2048x2_inst5_physical .INIT_0=256'b0010000001010100011000000001001000110000000100100110010000011110011101010011110000100000011110110100000000001011000000000101101001000001000110000000000000001011010100000010101101010000001010000001000001101110010100000010111000110000010111100111000000010110;
    SB_RAM40_4K \test_program.Ram2048x2_inst5_physical  (
            .RDATA({dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,instruction_11,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,instruction_10,dangling_wire_399,dangling_wire_400,dangling_wire_401}),
            .RADDR({N__12571,N__12733,N__12979,N__14170,N__13774,N__13987,N__13624,N__17674,N__15268,N__15658,N__15481}),
            .WADDR({N__12568,N__12730,N__12976,N__14161,N__13771,N__13978,N__13621,N__17671,N__15253,N__15655,N__15484}),
            .MASK({dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .WDATA({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .RCLKE(N__16221),
            .RCLK(N__33674),
            .RE(N__22555),
            .WCLKE(N__16220),
            .WCLK(N__33673),
            .WE());
    defparam \test_program.Ram2048x2_inst0_physical .WRITE_MODE=3;
    defparam \test_program.Ram2048x2_inst0_physical .READ_MODE=3;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_F=256'b0000100000101000000010000000000000000000000000000010011000100110000000110000000000000001000000110000001000010010000100110000000000110000001100010000000100100001001010000011101000111000001010000011101100111000001010010010101100001001000010000000101000101010;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_E=256'b0001111100011000000000000000011100101000001010000010001000000010000010100010010100000000000011100010000000100001001010100000111000001010001001010000000000001010000000000000000100011110000010100010001000100000000000000001000000110110001100100000001100000110;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_D=256'b0000011000000000000001010010010100000000000000110010000000100001000010000000101000011010000010100000110100001001000011010000100000011100000111000000110000001101000011010000100100100101001000000000110100100101000001000000000000001001000011010001000100101000;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_C=256'b0000111000001110000001000000000100001011000011110000001100000000000010010010111000000101000001000011101100001110000101110000010000001100000110100010100000101100000110100001101000111110000011000000110000011010001010000010110000101011001010110000111100011000;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_B=256'b0011100000101100001110000000101100001101000001010010011100111010001100010010010100001010000010100000111100000001000001010011111000011100000010000010101000001111000000110011000100000101000001100001110100011000000100110000111000000011000100000000000100000110;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_A=256'b0001100000011000001000100000011000001010000010000011010000000110000111000010100000000011001001110000100000001000001001110011111100101110000010000000100100101010000011000000100000101011001111100010101000001000000011010000111100011100000110000001101100001111;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_9=256'b0000101000010001000001000000111000010000000100010011101000001010000110100000010000110100001010000010010000001110000010000010100000000000000001000010110100111000001101100001111000110000000000010001111000110000000100000001100000111100001001000010000000000001;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_8=256'b0001100000100001000100000000000000001000000000000000000000000001000110000001000100000010000000100000110000010001000001110000111100011010000110000010110000001111000011000010110100001110000011100010111000101100001011010000111100001100001010000000101100001010;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_7=256'b0011111000000000000001000011101100000000000000010011101000111011001010100000000000000000001010000000000000001010000110000011100000010010000000100010000000110001001010100000101100000110001011000000010100000111001001000010010100001110000001100000011100000101;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_6=256'b0000110000000111000101010000010000001010000000110000001000000000000110000001001000000000001000000000101000010011001000100010000100101000000000110001000000110000000010110000001000110000001100010000100100100001000011100001111000101111001010010010110100001011;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_5=256'b0001100000111000000011110000111100101010001011000010110000001010000011000011100100001000000010010010110100100101001100110001101100000000001000000000111000011111001011110000010100000101001111100000110000001001000010110000100000010100000101000000100100001101;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_4=256'b0001010100001100000001010000000100000000000100000000010100000000000010000000100100011100000101000000010000001101000100000001000000001010000010000010100000011101000010000000000000000010000010000001000000110101000010000000100000101100001001000010110000000011;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_3=256'b0001000100110101000110000001100000100110001111100011010100010000000100000011111000010001000100000011001000110111001000000000010000011001001110000000001100011101000000100001001100110000001100010011101100010011000000100010001000011010000100110010000000110000;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_2=256'b0010101100000001000000010111000000011110011100110000101000101000000000010000100100001011000111000001001000010001000010000000000000000001000100110000000100011000011000100000001100100000001100000000000100100010000001000110101100010110001101000001100100001001;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_1=256'b0110100101110010001000100000110101000000011100100000100100001001001111010111011000100010000010110000000000000000010010010101100100011001001101100000100000001101001000100010011000101100010011000000000100101011000000010000011001101011011010000010000000000101;
    defparam \test_program.Ram2048x2_inst0_physical .INIT_0=256'b0000110001100011000100110000000000101100011001100011110100000001000000000010101001000010010101100000100000100000010101010000000100101000001001000010000001000000000011000011010000000011000000110111100001110010000110000000100001000000010110000000000000000010;
    SB_RAM40_4K \test_program.Ram2048x2_inst0_physical  (
            .RDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,instruction_1,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,instruction_0,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RADDR({N__12629,N__12791,N__13037,N__14225,N__13832,N__14042,N__13682,N__17732,N__15320,N__15716,N__15541}),
            .WADDR({N__12628,N__12790,N__13036,N__14221,N__13831,N__14038,N__13681,N__17731,N__15313,N__15715,N__15542}),
            .MASK({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463}),
            .WDATA({dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479}),
            .RCLKE(N__16233),
            .RCLK(N__33709),
            .RE(N__22479),
            .WCLKE(N__16232),
            .WCLK(N__33708),
            .WE());
    PRE_IO_GBUF CLK_3P3_MHZ_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__39684),
            .GLOBALBUFFEROUTPUT(CLK_3P3_MHZ_c_g));
    IO_PAD CLK_3P3_MHZ_ibuf_gb_io_iopad (
            .OE(N__39686),
            .DIN(N__39685),
            .DOUT(N__39684),
            .PACKAGEPIN(CLK_3P3_MHZ));
    defparam CLK_3P3_MHZ_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_3P3_MHZ_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_3P3_MHZ_ibuf_gb_io_preio (
            .PADOEN(N__39686),
            .PADOUT(N__39685),
            .PADIN(N__39684),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED1_obuf_iopad (
            .OE(N__39675),
            .DIN(N__39674),
            .DOUT(N__39673),
            .PACKAGEPIN(LED1));
    defparam LED1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED1_obuf_preio (
            .PADOEN(N__39675),
            .PADOUT(N__39674),
            .PADIN(N__39673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21032),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam BTN1_ibuf_iopad.PULLUP=1'b1;
    IO_PAD BTN1_ibuf_iopad (
            .OE(N__39666),
            .DIN(N__39665),
            .DOUT(N__39664),
            .PACKAGEPIN(BTN1));
    defparam BTN1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BTN1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BTN1_ibuf_preio (
            .PADOEN(N__39666),
            .PADOUT(N__39665),
            .PADIN(N__39664),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BTN1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__10148 (
            .O(N__39647),
            .I(N__39639));
    CascadeMux I__10147 (
            .O(N__39646),
            .I(N__39632));
    CascadeMux I__10146 (
            .O(N__39645),
            .I(N__39627));
    CascadeMux I__10145 (
            .O(N__39644),
            .I(N__39623));
    CascadeMux I__10144 (
            .O(N__39643),
            .I(N__39620));
    CascadeMux I__10143 (
            .O(N__39642),
            .I(N__39616));
    InMux I__10142 (
            .O(N__39639),
            .I(N__39613));
    CascadeMux I__10141 (
            .O(N__39638),
            .I(N__39610));
    InMux I__10140 (
            .O(N__39637),
            .I(N__39605));
    CascadeMux I__10139 (
            .O(N__39636),
            .I(N__39602));
    CascadeMux I__10138 (
            .O(N__39635),
            .I(N__39599));
    InMux I__10137 (
            .O(N__39632),
            .I(N__39588));
    InMux I__10136 (
            .O(N__39631),
            .I(N__39585));
    InMux I__10135 (
            .O(N__39630),
            .I(N__39582));
    InMux I__10134 (
            .O(N__39627),
            .I(N__39579));
    InMux I__10133 (
            .O(N__39626),
            .I(N__39576));
    InMux I__10132 (
            .O(N__39623),
            .I(N__39572));
    InMux I__10131 (
            .O(N__39620),
            .I(N__39569));
    CascadeMux I__10130 (
            .O(N__39619),
            .I(N__39565));
    InMux I__10129 (
            .O(N__39616),
            .I(N__39562));
    LocalMux I__10128 (
            .O(N__39613),
            .I(N__39559));
    InMux I__10127 (
            .O(N__39610),
            .I(N__39556));
    InMux I__10126 (
            .O(N__39609),
            .I(N__39553));
    InMux I__10125 (
            .O(N__39608),
            .I(N__39550));
    LocalMux I__10124 (
            .O(N__39605),
            .I(N__39547));
    InMux I__10123 (
            .O(N__39602),
            .I(N__39539));
    InMux I__10122 (
            .O(N__39599),
            .I(N__39536));
    CascadeMux I__10121 (
            .O(N__39598),
            .I(N__39532));
    CascadeMux I__10120 (
            .O(N__39597),
            .I(N__39529));
    InMux I__10119 (
            .O(N__39596),
            .I(N__39526));
    InMux I__10118 (
            .O(N__39595),
            .I(N__39523));
    CascadeMux I__10117 (
            .O(N__39594),
            .I(N__39520));
    CascadeMux I__10116 (
            .O(N__39593),
            .I(N__39517));
    InMux I__10115 (
            .O(N__39592),
            .I(N__39514));
    InMux I__10114 (
            .O(N__39591),
            .I(N__39511));
    LocalMux I__10113 (
            .O(N__39588),
            .I(N__39508));
    LocalMux I__10112 (
            .O(N__39585),
            .I(N__39503));
    LocalMux I__10111 (
            .O(N__39582),
            .I(N__39503));
    LocalMux I__10110 (
            .O(N__39579),
            .I(N__39498));
    LocalMux I__10109 (
            .O(N__39576),
            .I(N__39498));
    CascadeMux I__10108 (
            .O(N__39575),
            .I(N__39495));
    LocalMux I__10107 (
            .O(N__39572),
            .I(N__39489));
    LocalMux I__10106 (
            .O(N__39569),
            .I(N__39489));
    InMux I__10105 (
            .O(N__39568),
            .I(N__39486));
    InMux I__10104 (
            .O(N__39565),
            .I(N__39483));
    LocalMux I__10103 (
            .O(N__39562),
            .I(N__39478));
    Span4Mux_v I__10102 (
            .O(N__39559),
            .I(N__39478));
    LocalMux I__10101 (
            .O(N__39556),
            .I(N__39469));
    LocalMux I__10100 (
            .O(N__39553),
            .I(N__39469));
    LocalMux I__10099 (
            .O(N__39550),
            .I(N__39469));
    Span4Mux_v I__10098 (
            .O(N__39547),
            .I(N__39469));
    CascadeMux I__10097 (
            .O(N__39546),
            .I(N__39466));
    InMux I__10096 (
            .O(N__39545),
            .I(N__39463));
    InMux I__10095 (
            .O(N__39544),
            .I(N__39460));
    CascadeMux I__10094 (
            .O(N__39543),
            .I(N__39457));
    CascadeMux I__10093 (
            .O(N__39542),
            .I(N__39454));
    LocalMux I__10092 (
            .O(N__39539),
            .I(N__39451));
    LocalMux I__10091 (
            .O(N__39536),
            .I(N__39447));
    InMux I__10090 (
            .O(N__39535),
            .I(N__39444));
    InMux I__10089 (
            .O(N__39532),
            .I(N__39441));
    InMux I__10088 (
            .O(N__39529),
            .I(N__39438));
    LocalMux I__10087 (
            .O(N__39526),
            .I(N__39435));
    LocalMux I__10086 (
            .O(N__39523),
            .I(N__39432));
    InMux I__10085 (
            .O(N__39520),
            .I(N__39429));
    InMux I__10084 (
            .O(N__39517),
            .I(N__39426));
    LocalMux I__10083 (
            .O(N__39514),
            .I(N__39423));
    LocalMux I__10082 (
            .O(N__39511),
            .I(N__39416));
    Span4Mux_s3_h I__10081 (
            .O(N__39508),
            .I(N__39416));
    Span4Mux_v I__10080 (
            .O(N__39503),
            .I(N__39416));
    Span4Mux_s3_v I__10079 (
            .O(N__39498),
            .I(N__39413));
    InMux I__10078 (
            .O(N__39495),
            .I(N__39410));
    InMux I__10077 (
            .O(N__39494),
            .I(N__39407));
    Span4Mux_s3_v I__10076 (
            .O(N__39489),
            .I(N__39402));
    LocalMux I__10075 (
            .O(N__39486),
            .I(N__39402));
    LocalMux I__10074 (
            .O(N__39483),
            .I(N__39395));
    Span4Mux_s0_h I__10073 (
            .O(N__39478),
            .I(N__39395));
    Span4Mux_v I__10072 (
            .O(N__39469),
            .I(N__39395));
    InMux I__10071 (
            .O(N__39466),
            .I(N__39392));
    LocalMux I__10070 (
            .O(N__39463),
            .I(N__39389));
    LocalMux I__10069 (
            .O(N__39460),
            .I(N__39386));
    InMux I__10068 (
            .O(N__39457),
            .I(N__39383));
    InMux I__10067 (
            .O(N__39454),
            .I(N__39380));
    Span4Mux_v I__10066 (
            .O(N__39451),
            .I(N__39377));
    InMux I__10065 (
            .O(N__39450),
            .I(N__39374));
    Sp12to4 I__10064 (
            .O(N__39447),
            .I(N__39369));
    LocalMux I__10063 (
            .O(N__39444),
            .I(N__39369));
    LocalMux I__10062 (
            .O(N__39441),
            .I(N__39366));
    LocalMux I__10061 (
            .O(N__39438),
            .I(N__39359));
    Span4Mux_v I__10060 (
            .O(N__39435),
            .I(N__39359));
    Span4Mux_h I__10059 (
            .O(N__39432),
            .I(N__39359));
    LocalMux I__10058 (
            .O(N__39429),
            .I(N__39350));
    LocalMux I__10057 (
            .O(N__39426),
            .I(N__39350));
    Span4Mux_h I__10056 (
            .O(N__39423),
            .I(N__39350));
    Span4Mux_h I__10055 (
            .O(N__39416),
            .I(N__39350));
    Span4Mux_h I__10054 (
            .O(N__39413),
            .I(N__39345));
    LocalMux I__10053 (
            .O(N__39410),
            .I(N__39345));
    LocalMux I__10052 (
            .O(N__39407),
            .I(N__39342));
    Span4Mux_v I__10051 (
            .O(N__39402),
            .I(N__39335));
    Span4Mux_h I__10050 (
            .O(N__39395),
            .I(N__39335));
    LocalMux I__10049 (
            .O(N__39392),
            .I(N__39335));
    Span4Mux_v I__10048 (
            .O(N__39389),
            .I(N__39330));
    Span4Mux_v I__10047 (
            .O(N__39386),
            .I(N__39330));
    LocalMux I__10046 (
            .O(N__39383),
            .I(N__39321));
    LocalMux I__10045 (
            .O(N__39380),
            .I(N__39321));
    Sp12to4 I__10044 (
            .O(N__39377),
            .I(N__39321));
    LocalMux I__10043 (
            .O(N__39374),
            .I(N__39321));
    Span12Mux_s5_v I__10042 (
            .O(N__39369),
            .I(N__39318));
    Span4Mux_s3_h I__10041 (
            .O(N__39366),
            .I(N__39313));
    Span4Mux_h I__10040 (
            .O(N__39359),
            .I(N__39313));
    Span4Mux_v I__10039 (
            .O(N__39350),
            .I(N__39308));
    Span4Mux_s3_v I__10038 (
            .O(N__39345),
            .I(N__39308));
    Span4Mux_h I__10037 (
            .O(N__39342),
            .I(N__39303));
    Span4Mux_h I__10036 (
            .O(N__39335),
            .I(N__39303));
    Odrv4 I__10035 (
            .O(N__39330),
            .I(\processor_zipi8.arith_logical_result_1 ));
    Odrv12 I__10034 (
            .O(N__39321),
            .I(\processor_zipi8.arith_logical_result_1 ));
    Odrv12 I__10033 (
            .O(N__39318),
            .I(\processor_zipi8.arith_logical_result_1 ));
    Odrv4 I__10032 (
            .O(N__39313),
            .I(\processor_zipi8.arith_logical_result_1 ));
    Odrv4 I__10031 (
            .O(N__39308),
            .I(\processor_zipi8.arith_logical_result_1 ));
    Odrv4 I__10030 (
            .O(N__39303),
            .I(\processor_zipi8.arith_logical_result_1 ));
    CascadeMux I__10029 (
            .O(N__39290),
            .I(N__39286));
    CascadeMux I__10028 (
            .O(N__39289),
            .I(N__39279));
    InMux I__10027 (
            .O(N__39286),
            .I(N__39276));
    CascadeMux I__10026 (
            .O(N__39285),
            .I(N__39273));
    CascadeMux I__10025 (
            .O(N__39284),
            .I(N__39270));
    CascadeMux I__10024 (
            .O(N__39283),
            .I(N__39267));
    CascadeMux I__10023 (
            .O(N__39282),
            .I(N__39264));
    InMux I__10022 (
            .O(N__39279),
            .I(N__39255));
    LocalMux I__10021 (
            .O(N__39276),
            .I(N__39252));
    InMux I__10020 (
            .O(N__39273),
            .I(N__39249));
    InMux I__10019 (
            .O(N__39270),
            .I(N__39244));
    InMux I__10018 (
            .O(N__39267),
            .I(N__39237));
    InMux I__10017 (
            .O(N__39264),
            .I(N__39234));
    InMux I__10016 (
            .O(N__39263),
            .I(N__39230));
    CascadeMux I__10015 (
            .O(N__39262),
            .I(N__39221));
    InMux I__10014 (
            .O(N__39261),
            .I(N__39218));
    CascadeMux I__10013 (
            .O(N__39260),
            .I(N__39215));
    InMux I__10012 (
            .O(N__39259),
            .I(N__39212));
    InMux I__10011 (
            .O(N__39258),
            .I(N__39209));
    LocalMux I__10010 (
            .O(N__39255),
            .I(N__39202));
    Span4Mux_h I__10009 (
            .O(N__39252),
            .I(N__39202));
    LocalMux I__10008 (
            .O(N__39249),
            .I(N__39202));
    CascadeMux I__10007 (
            .O(N__39248),
            .I(N__39199));
    InMux I__10006 (
            .O(N__39247),
            .I(N__39195));
    LocalMux I__10005 (
            .O(N__39244),
            .I(N__39192));
    InMux I__10004 (
            .O(N__39243),
            .I(N__39189));
    InMux I__10003 (
            .O(N__39242),
            .I(N__39185));
    InMux I__10002 (
            .O(N__39241),
            .I(N__39182));
    InMux I__10001 (
            .O(N__39240),
            .I(N__39179));
    LocalMux I__10000 (
            .O(N__39237),
            .I(N__39172));
    LocalMux I__9999 (
            .O(N__39234),
            .I(N__39172));
    CascadeMux I__9998 (
            .O(N__39233),
            .I(N__39169));
    LocalMux I__9997 (
            .O(N__39230),
            .I(N__39166));
    CascadeMux I__9996 (
            .O(N__39229),
            .I(N__39163));
    CascadeMux I__9995 (
            .O(N__39228),
            .I(N__39160));
    CascadeMux I__9994 (
            .O(N__39227),
            .I(N__39157));
    InMux I__9993 (
            .O(N__39226),
            .I(N__39154));
    InMux I__9992 (
            .O(N__39225),
            .I(N__39151));
    InMux I__9991 (
            .O(N__39224),
            .I(N__39148));
    InMux I__9990 (
            .O(N__39221),
            .I(N__39145));
    LocalMux I__9989 (
            .O(N__39218),
            .I(N__39142));
    InMux I__9988 (
            .O(N__39215),
            .I(N__39139));
    LocalMux I__9987 (
            .O(N__39212),
            .I(N__39136));
    LocalMux I__9986 (
            .O(N__39209),
            .I(N__39131));
    Span4Mux_s2_h I__9985 (
            .O(N__39202),
            .I(N__39131));
    InMux I__9984 (
            .O(N__39199),
            .I(N__39128));
    InMux I__9983 (
            .O(N__39198),
            .I(N__39124));
    LocalMux I__9982 (
            .O(N__39195),
            .I(N__39121));
    Span4Mux_v I__9981 (
            .O(N__39192),
            .I(N__39116));
    LocalMux I__9980 (
            .O(N__39189),
            .I(N__39116));
    InMux I__9979 (
            .O(N__39188),
            .I(N__39113));
    LocalMux I__9978 (
            .O(N__39185),
            .I(N__39110));
    LocalMux I__9977 (
            .O(N__39182),
            .I(N__39107));
    LocalMux I__9976 (
            .O(N__39179),
            .I(N__39104));
    InMux I__9975 (
            .O(N__39178),
            .I(N__39101));
    InMux I__9974 (
            .O(N__39177),
            .I(N__39098));
    Span4Mux_h I__9973 (
            .O(N__39172),
            .I(N__39095));
    InMux I__9972 (
            .O(N__39169),
            .I(N__39091));
    IoSpan4Mux I__9971 (
            .O(N__39166),
            .I(N__39088));
    InMux I__9970 (
            .O(N__39163),
            .I(N__39085));
    InMux I__9969 (
            .O(N__39160),
            .I(N__39082));
    InMux I__9968 (
            .O(N__39157),
            .I(N__39079));
    LocalMux I__9967 (
            .O(N__39154),
            .I(N__39074));
    LocalMux I__9966 (
            .O(N__39151),
            .I(N__39074));
    LocalMux I__9965 (
            .O(N__39148),
            .I(N__39071));
    LocalMux I__9964 (
            .O(N__39145),
            .I(N__39068));
    Span4Mux_s2_h I__9963 (
            .O(N__39142),
            .I(N__39059));
    LocalMux I__9962 (
            .O(N__39139),
            .I(N__39059));
    Span4Mux_s2_h I__9961 (
            .O(N__39136),
            .I(N__39059));
    Span4Mux_v I__9960 (
            .O(N__39131),
            .I(N__39059));
    LocalMux I__9959 (
            .O(N__39128),
            .I(N__39056));
    InMux I__9958 (
            .O(N__39127),
            .I(N__39053));
    LocalMux I__9957 (
            .O(N__39124),
            .I(N__39049));
    Span4Mux_h I__9956 (
            .O(N__39121),
            .I(N__39044));
    Span4Mux_s1_h I__9955 (
            .O(N__39116),
            .I(N__39044));
    LocalMux I__9954 (
            .O(N__39113),
            .I(N__39039));
    Span4Mux_s1_h I__9953 (
            .O(N__39110),
            .I(N__39039));
    Span4Mux_h I__9952 (
            .O(N__39107),
            .I(N__39032));
    Span4Mux_h I__9951 (
            .O(N__39104),
            .I(N__39032));
    LocalMux I__9950 (
            .O(N__39101),
            .I(N__39032));
    LocalMux I__9949 (
            .O(N__39098),
            .I(N__39029));
    Sp12to4 I__9948 (
            .O(N__39095),
            .I(N__39026));
    InMux I__9947 (
            .O(N__39094),
            .I(N__39023));
    LocalMux I__9946 (
            .O(N__39091),
            .I(N__39020));
    Span4Mux_s2_h I__9945 (
            .O(N__39088),
            .I(N__39015));
    LocalMux I__9944 (
            .O(N__39085),
            .I(N__39015));
    LocalMux I__9943 (
            .O(N__39082),
            .I(N__39012));
    LocalMux I__9942 (
            .O(N__39079),
            .I(N__39007));
    Span4Mux_h I__9941 (
            .O(N__39074),
            .I(N__39007));
    Span4Mux_h I__9940 (
            .O(N__39071),
            .I(N__39000));
    Span4Mux_v I__9939 (
            .O(N__39068),
            .I(N__39000));
    Span4Mux_h I__9938 (
            .O(N__39059),
            .I(N__39000));
    Span4Mux_h I__9937 (
            .O(N__39056),
            .I(N__38995));
    LocalMux I__9936 (
            .O(N__39053),
            .I(N__38995));
    InMux I__9935 (
            .O(N__39052),
            .I(N__38992));
    Span12Mux_s6_h I__9934 (
            .O(N__39049),
            .I(N__38989));
    Span4Mux_h I__9933 (
            .O(N__39044),
            .I(N__38982));
    Span4Mux_h I__9932 (
            .O(N__39039),
            .I(N__38982));
    Span4Mux_v I__9931 (
            .O(N__39032),
            .I(N__38982));
    Span12Mux_s1_h I__9930 (
            .O(N__39029),
            .I(N__38977));
    Span12Mux_s8_v I__9929 (
            .O(N__39026),
            .I(N__38977));
    LocalMux I__9928 (
            .O(N__39023),
            .I(N__38970));
    Span4Mux_h I__9927 (
            .O(N__39020),
            .I(N__38970));
    Span4Mux_h I__9926 (
            .O(N__39015),
            .I(N__38970));
    Span12Mux_s5_h I__9925 (
            .O(N__39012),
            .I(N__38961));
    Sp12to4 I__9924 (
            .O(N__39007),
            .I(N__38961));
    Sp12to4 I__9923 (
            .O(N__39000),
            .I(N__38961));
    Sp12to4 I__9922 (
            .O(N__38995),
            .I(N__38961));
    LocalMux I__9921 (
            .O(N__38992),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ));
    Odrv12 I__9920 (
            .O(N__38989),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ));
    Odrv4 I__9919 (
            .O(N__38982),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ));
    Odrv12 I__9918 (
            .O(N__38977),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ));
    Odrv4 I__9917 (
            .O(N__38970),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ));
    Odrv12 I__9916 (
            .O(N__38961),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ));
    CascadeMux I__9915 (
            .O(N__38948),
            .I(N__38945));
    InMux I__9914 (
            .O(N__38945),
            .I(N__38942));
    LocalMux I__9913 (
            .O(N__38942),
            .I(N__38938));
    InMux I__9912 (
            .O(N__38941),
            .I(N__38935));
    Span4Mux_v I__9911 (
            .O(N__38938),
            .I(N__38932));
    LocalMux I__9910 (
            .O(N__38935),
            .I(N__38929));
    Odrv4 I__9909 (
            .O(N__38932),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1 ));
    Odrv12 I__9908 (
            .O(N__38929),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1 ));
    InMux I__9907 (
            .O(N__38924),
            .I(N__38921));
    LocalMux I__9906 (
            .O(N__38921),
            .I(N__38917));
    InMux I__9905 (
            .O(N__38920),
            .I(N__38914));
    Odrv4 I__9904 (
            .O(N__38917),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1 ));
    LocalMux I__9903 (
            .O(N__38914),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1 ));
    CascadeMux I__9902 (
            .O(N__38909),
            .I(N__38906));
    InMux I__9901 (
            .O(N__38906),
            .I(N__38903));
    LocalMux I__9900 (
            .O(N__38903),
            .I(N__38900));
    Span4Mux_h I__9899 (
            .O(N__38900),
            .I(N__38897));
    Span4Mux_s0_h I__9898 (
            .O(N__38897),
            .I(N__38894));
    Odrv4 I__9897 (
            .O(N__38894),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_1 ));
    CascadeMux I__9896 (
            .O(N__38891),
            .I(N__38883));
    CascadeMux I__9895 (
            .O(N__38890),
            .I(N__38875));
    InMux I__9894 (
            .O(N__38889),
            .I(N__38871));
    CascadeMux I__9893 (
            .O(N__38888),
            .I(N__38868));
    InMux I__9892 (
            .O(N__38887),
            .I(N__38864));
    InMux I__9891 (
            .O(N__38886),
            .I(N__38861));
    InMux I__9890 (
            .O(N__38883),
            .I(N__38858));
    InMux I__9889 (
            .O(N__38882),
            .I(N__38855));
    CascadeMux I__9888 (
            .O(N__38881),
            .I(N__38852));
    CascadeMux I__9887 (
            .O(N__38880),
            .I(N__38848));
    CascadeMux I__9886 (
            .O(N__38879),
            .I(N__38844));
    InMux I__9885 (
            .O(N__38878),
            .I(N__38840));
    InMux I__9884 (
            .O(N__38875),
            .I(N__38837));
    InMux I__9883 (
            .O(N__38874),
            .I(N__38827));
    LocalMux I__9882 (
            .O(N__38871),
            .I(N__38824));
    InMux I__9881 (
            .O(N__38868),
            .I(N__38821));
    InMux I__9880 (
            .O(N__38867),
            .I(N__38817));
    LocalMux I__9879 (
            .O(N__38864),
            .I(N__38814));
    LocalMux I__9878 (
            .O(N__38861),
            .I(N__38811));
    LocalMux I__9877 (
            .O(N__38858),
            .I(N__38806));
    LocalMux I__9876 (
            .O(N__38855),
            .I(N__38806));
    InMux I__9875 (
            .O(N__38852),
            .I(N__38803));
    InMux I__9874 (
            .O(N__38851),
            .I(N__38796));
    InMux I__9873 (
            .O(N__38848),
            .I(N__38793));
    InMux I__9872 (
            .O(N__38847),
            .I(N__38790));
    InMux I__9871 (
            .O(N__38844),
            .I(N__38787));
    CascadeMux I__9870 (
            .O(N__38843),
            .I(N__38784));
    LocalMux I__9869 (
            .O(N__38840),
            .I(N__38779));
    LocalMux I__9868 (
            .O(N__38837),
            .I(N__38776));
    InMux I__9867 (
            .O(N__38836),
            .I(N__38773));
    InMux I__9866 (
            .O(N__38835),
            .I(N__38770));
    InMux I__9865 (
            .O(N__38834),
            .I(N__38767));
    CascadeMux I__9864 (
            .O(N__38833),
            .I(N__38764));
    InMux I__9863 (
            .O(N__38832),
            .I(N__38761));
    InMux I__9862 (
            .O(N__38831),
            .I(N__38758));
    InMux I__9861 (
            .O(N__38830),
            .I(N__38755));
    LocalMux I__9860 (
            .O(N__38827),
            .I(N__38752));
    Span4Mux_v I__9859 (
            .O(N__38824),
            .I(N__38747));
    LocalMux I__9858 (
            .O(N__38821),
            .I(N__38747));
    InMux I__9857 (
            .O(N__38820),
            .I(N__38744));
    LocalMux I__9856 (
            .O(N__38817),
            .I(N__38739));
    Span4Mux_s3_h I__9855 (
            .O(N__38814),
            .I(N__38739));
    Span4Mux_v I__9854 (
            .O(N__38811),
            .I(N__38732));
    Span4Mux_s3_h I__9853 (
            .O(N__38806),
            .I(N__38732));
    LocalMux I__9852 (
            .O(N__38803),
            .I(N__38732));
    CascadeMux I__9851 (
            .O(N__38802),
            .I(N__38726));
    InMux I__9850 (
            .O(N__38801),
            .I(N__38722));
    InMux I__9849 (
            .O(N__38800),
            .I(N__38719));
    InMux I__9848 (
            .O(N__38799),
            .I(N__38716));
    LocalMux I__9847 (
            .O(N__38796),
            .I(N__38711));
    LocalMux I__9846 (
            .O(N__38793),
            .I(N__38711));
    LocalMux I__9845 (
            .O(N__38790),
            .I(N__38706));
    LocalMux I__9844 (
            .O(N__38787),
            .I(N__38706));
    InMux I__9843 (
            .O(N__38784),
            .I(N__38703));
    InMux I__9842 (
            .O(N__38783),
            .I(N__38700));
    InMux I__9841 (
            .O(N__38782),
            .I(N__38697));
    Span4Mux_h I__9840 (
            .O(N__38779),
            .I(N__38686));
    Span4Mux_s3_h I__9839 (
            .O(N__38776),
            .I(N__38686));
    LocalMux I__9838 (
            .O(N__38773),
            .I(N__38686));
    LocalMux I__9837 (
            .O(N__38770),
            .I(N__38686));
    LocalMux I__9836 (
            .O(N__38767),
            .I(N__38686));
    InMux I__9835 (
            .O(N__38764),
            .I(N__38683));
    LocalMux I__9834 (
            .O(N__38761),
            .I(N__38678));
    LocalMux I__9833 (
            .O(N__38758),
            .I(N__38678));
    LocalMux I__9832 (
            .O(N__38755),
            .I(N__38673));
    Span4Mux_s2_v I__9831 (
            .O(N__38752),
            .I(N__38673));
    Span4Mux_s1_h I__9830 (
            .O(N__38747),
            .I(N__38670));
    LocalMux I__9829 (
            .O(N__38744),
            .I(N__38663));
    Span4Mux_v I__9828 (
            .O(N__38739),
            .I(N__38663));
    Span4Mux_h I__9827 (
            .O(N__38732),
            .I(N__38663));
    CascadeMux I__9826 (
            .O(N__38731),
            .I(N__38660));
    InMux I__9825 (
            .O(N__38730),
            .I(N__38657));
    InMux I__9824 (
            .O(N__38729),
            .I(N__38654));
    InMux I__9823 (
            .O(N__38726),
            .I(N__38651));
    InMux I__9822 (
            .O(N__38725),
            .I(N__38648));
    LocalMux I__9821 (
            .O(N__38722),
            .I(N__38641));
    LocalMux I__9820 (
            .O(N__38719),
            .I(N__38641));
    LocalMux I__9819 (
            .O(N__38716),
            .I(N__38641));
    Span4Mux_v I__9818 (
            .O(N__38711),
            .I(N__38636));
    Span4Mux_s2_v I__9817 (
            .O(N__38706),
            .I(N__38636));
    LocalMux I__9816 (
            .O(N__38703),
            .I(N__38633));
    LocalMux I__9815 (
            .O(N__38700),
            .I(N__38626));
    LocalMux I__9814 (
            .O(N__38697),
            .I(N__38626));
    Sp12to4 I__9813 (
            .O(N__38686),
            .I(N__38626));
    LocalMux I__9812 (
            .O(N__38683),
            .I(N__38617));
    Span4Mux_v I__9811 (
            .O(N__38678),
            .I(N__38617));
    Span4Mux_v I__9810 (
            .O(N__38673),
            .I(N__38617));
    Span4Mux_v I__9809 (
            .O(N__38670),
            .I(N__38617));
    Sp12to4 I__9808 (
            .O(N__38663),
            .I(N__38614));
    InMux I__9807 (
            .O(N__38660),
            .I(N__38611));
    LocalMux I__9806 (
            .O(N__38657),
            .I(N__38604));
    LocalMux I__9805 (
            .O(N__38654),
            .I(N__38604));
    LocalMux I__9804 (
            .O(N__38651),
            .I(N__38604));
    LocalMux I__9803 (
            .O(N__38648),
            .I(N__38599));
    Span12Mux_s10_h I__9802 (
            .O(N__38641),
            .I(N__38599));
    Span4Mux_v I__9801 (
            .O(N__38636),
            .I(N__38596));
    Span12Mux_s3_h I__9800 (
            .O(N__38633),
            .I(N__38585));
    Span12Mux_s6_v I__9799 (
            .O(N__38626),
            .I(N__38585));
    Sp12to4 I__9798 (
            .O(N__38617),
            .I(N__38585));
    Span12Mux_s9_v I__9797 (
            .O(N__38614),
            .I(N__38585));
    LocalMux I__9796 (
            .O(N__38611),
            .I(N__38585));
    Odrv12 I__9795 (
            .O(N__38604),
            .I(\processor_zipi8.arith_logical_result_2 ));
    Odrv12 I__9794 (
            .O(N__38599),
            .I(\processor_zipi8.arith_logical_result_2 ));
    Odrv4 I__9793 (
            .O(N__38596),
            .I(\processor_zipi8.arith_logical_result_2 ));
    Odrv12 I__9792 (
            .O(N__38585),
            .I(\processor_zipi8.arith_logical_result_2 ));
    CascadeMux I__9791 (
            .O(N__38576),
            .I(N__38571));
    InMux I__9790 (
            .O(N__38575),
            .I(N__38562));
    InMux I__9789 (
            .O(N__38574),
            .I(N__38559));
    InMux I__9788 (
            .O(N__38571),
            .I(N__38553));
    CascadeMux I__9787 (
            .O(N__38570),
            .I(N__38546));
    CascadeMux I__9786 (
            .O(N__38569),
            .I(N__38542));
    CascadeMux I__9785 (
            .O(N__38568),
            .I(N__38537));
    CascadeMux I__9784 (
            .O(N__38567),
            .I(N__38534));
    InMux I__9783 (
            .O(N__38566),
            .I(N__38527));
    InMux I__9782 (
            .O(N__38565),
            .I(N__38524));
    LocalMux I__9781 (
            .O(N__38562),
            .I(N__38519));
    LocalMux I__9780 (
            .O(N__38559),
            .I(N__38519));
    CascadeMux I__9779 (
            .O(N__38558),
            .I(N__38514));
    InMux I__9778 (
            .O(N__38557),
            .I(N__38510));
    InMux I__9777 (
            .O(N__38556),
            .I(N__38507));
    LocalMux I__9776 (
            .O(N__38553),
            .I(N__38502));
    CascadeMux I__9775 (
            .O(N__38552),
            .I(N__38499));
    InMux I__9774 (
            .O(N__38551),
            .I(N__38496));
    InMux I__9773 (
            .O(N__38550),
            .I(N__38493));
    InMux I__9772 (
            .O(N__38549),
            .I(N__38490));
    InMux I__9771 (
            .O(N__38546),
            .I(N__38487));
    InMux I__9770 (
            .O(N__38545),
            .I(N__38484));
    InMux I__9769 (
            .O(N__38542),
            .I(N__38481));
    InMux I__9768 (
            .O(N__38541),
            .I(N__38478));
    CascadeMux I__9767 (
            .O(N__38540),
            .I(N__38475));
    InMux I__9766 (
            .O(N__38537),
            .I(N__38472));
    InMux I__9765 (
            .O(N__38534),
            .I(N__38469));
    InMux I__9764 (
            .O(N__38533),
            .I(N__38466));
    CascadeMux I__9763 (
            .O(N__38532),
            .I(N__38463));
    CascadeMux I__9762 (
            .O(N__38531),
            .I(N__38458));
    CascadeMux I__9761 (
            .O(N__38530),
            .I(N__38455));
    LocalMux I__9760 (
            .O(N__38527),
            .I(N__38452));
    LocalMux I__9759 (
            .O(N__38524),
            .I(N__38447));
    Span4Mux_v I__9758 (
            .O(N__38519),
            .I(N__38447));
    CascadeMux I__9757 (
            .O(N__38518),
            .I(N__38443));
    CascadeMux I__9756 (
            .O(N__38517),
            .I(N__38440));
    InMux I__9755 (
            .O(N__38514),
            .I(N__38437));
    InMux I__9754 (
            .O(N__38513),
            .I(N__38434));
    LocalMux I__9753 (
            .O(N__38510),
            .I(N__38429));
    LocalMux I__9752 (
            .O(N__38507),
            .I(N__38429));
    CascadeMux I__9751 (
            .O(N__38506),
            .I(N__38426));
    InMux I__9750 (
            .O(N__38505),
            .I(N__38422));
    Span4Mux_v I__9749 (
            .O(N__38502),
            .I(N__38419));
    InMux I__9748 (
            .O(N__38499),
            .I(N__38416));
    LocalMux I__9747 (
            .O(N__38496),
            .I(N__38411));
    LocalMux I__9746 (
            .O(N__38493),
            .I(N__38411));
    LocalMux I__9745 (
            .O(N__38490),
            .I(N__38406));
    LocalMux I__9744 (
            .O(N__38487),
            .I(N__38406));
    LocalMux I__9743 (
            .O(N__38484),
            .I(N__38403));
    LocalMux I__9742 (
            .O(N__38481),
            .I(N__38398));
    LocalMux I__9741 (
            .O(N__38478),
            .I(N__38398));
    InMux I__9740 (
            .O(N__38475),
            .I(N__38395));
    LocalMux I__9739 (
            .O(N__38472),
            .I(N__38388));
    LocalMux I__9738 (
            .O(N__38469),
            .I(N__38388));
    LocalMux I__9737 (
            .O(N__38466),
            .I(N__38388));
    InMux I__9736 (
            .O(N__38463),
            .I(N__38385));
    InMux I__9735 (
            .O(N__38462),
            .I(N__38382));
    CascadeMux I__9734 (
            .O(N__38461),
            .I(N__38379));
    InMux I__9733 (
            .O(N__38458),
            .I(N__38376));
    InMux I__9732 (
            .O(N__38455),
            .I(N__38373));
    Span4Mux_v I__9731 (
            .O(N__38452),
            .I(N__38368));
    Span4Mux_v I__9730 (
            .O(N__38447),
            .I(N__38368));
    InMux I__9729 (
            .O(N__38446),
            .I(N__38365));
    InMux I__9728 (
            .O(N__38443),
            .I(N__38362));
    InMux I__9727 (
            .O(N__38440),
            .I(N__38359));
    LocalMux I__9726 (
            .O(N__38437),
            .I(N__38352));
    LocalMux I__9725 (
            .O(N__38434),
            .I(N__38352));
    Span4Mux_v I__9724 (
            .O(N__38429),
            .I(N__38352));
    InMux I__9723 (
            .O(N__38426),
            .I(N__38349));
    InMux I__9722 (
            .O(N__38425),
            .I(N__38346));
    LocalMux I__9721 (
            .O(N__38422),
            .I(N__38341));
    Span4Mux_v I__9720 (
            .O(N__38419),
            .I(N__38341));
    LocalMux I__9719 (
            .O(N__38416),
            .I(N__38334));
    Span4Mux_v I__9718 (
            .O(N__38411),
            .I(N__38334));
    Span4Mux_s3_h I__9717 (
            .O(N__38406),
            .I(N__38334));
    Span4Mux_v I__9716 (
            .O(N__38403),
            .I(N__38325));
    Span4Mux_s3_h I__9715 (
            .O(N__38398),
            .I(N__38325));
    LocalMux I__9714 (
            .O(N__38395),
            .I(N__38325));
    Span4Mux_v I__9713 (
            .O(N__38388),
            .I(N__38325));
    LocalMux I__9712 (
            .O(N__38385),
            .I(N__38320));
    LocalMux I__9711 (
            .O(N__38382),
            .I(N__38320));
    InMux I__9710 (
            .O(N__38379),
            .I(N__38317));
    LocalMux I__9709 (
            .O(N__38376),
            .I(N__38314));
    LocalMux I__9708 (
            .O(N__38373),
            .I(N__38311));
    Span4Mux_h I__9707 (
            .O(N__38368),
            .I(N__38307));
    LocalMux I__9706 (
            .O(N__38365),
            .I(N__38302));
    LocalMux I__9705 (
            .O(N__38362),
            .I(N__38302));
    LocalMux I__9704 (
            .O(N__38359),
            .I(N__38299));
    Span4Mux_v I__9703 (
            .O(N__38352),
            .I(N__38296));
    LocalMux I__9702 (
            .O(N__38349),
            .I(N__38289));
    LocalMux I__9701 (
            .O(N__38346),
            .I(N__38289));
    Span4Mux_v I__9700 (
            .O(N__38341),
            .I(N__38289));
    Span4Mux_h I__9699 (
            .O(N__38334),
            .I(N__38282));
    Span4Mux_h I__9698 (
            .O(N__38325),
            .I(N__38282));
    Span4Mux_v I__9697 (
            .O(N__38320),
            .I(N__38282));
    LocalMux I__9696 (
            .O(N__38317),
            .I(N__38279));
    Span4Mux_s3_v I__9695 (
            .O(N__38314),
            .I(N__38274));
    Span4Mux_v I__9694 (
            .O(N__38311),
            .I(N__38274));
    InMux I__9693 (
            .O(N__38310),
            .I(N__38271));
    Span4Mux_h I__9692 (
            .O(N__38307),
            .I(N__38268));
    Span4Mux_s2_v I__9691 (
            .O(N__38302),
            .I(N__38259));
    Span4Mux_h I__9690 (
            .O(N__38299),
            .I(N__38259));
    Span4Mux_v I__9689 (
            .O(N__38296),
            .I(N__38259));
    Span4Mux_h I__9688 (
            .O(N__38289),
            .I(N__38259));
    Span4Mux_v I__9687 (
            .O(N__38282),
            .I(N__38256));
    Span4Mux_h I__9686 (
            .O(N__38279),
            .I(N__38249));
    Span4Mux_h I__9685 (
            .O(N__38274),
            .I(N__38249));
    LocalMux I__9684 (
            .O(N__38271),
            .I(N__38249));
    Odrv4 I__9683 (
            .O(N__38268),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265 ));
    Odrv4 I__9682 (
            .O(N__38259),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265 ));
    Odrv4 I__9681 (
            .O(N__38256),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265 ));
    Odrv4 I__9680 (
            .O(N__38249),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265 ));
    InMux I__9679 (
            .O(N__38240),
            .I(N__38237));
    LocalMux I__9678 (
            .O(N__38237),
            .I(N__38233));
    InMux I__9677 (
            .O(N__38236),
            .I(N__38230));
    Span4Mux_s3_h I__9676 (
            .O(N__38233),
            .I(N__38227));
    LocalMux I__9675 (
            .O(N__38230),
            .I(N__38224));
    Odrv4 I__9674 (
            .O(N__38227),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2 ));
    Odrv12 I__9673 (
            .O(N__38224),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2 ));
    InMux I__9672 (
            .O(N__38219),
            .I(N__38216));
    LocalMux I__9671 (
            .O(N__38216),
            .I(N__38212));
    InMux I__9670 (
            .O(N__38215),
            .I(N__38209));
    Odrv4 I__9669 (
            .O(N__38212),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2 ));
    LocalMux I__9668 (
            .O(N__38209),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2 ));
    InMux I__9667 (
            .O(N__38204),
            .I(N__38201));
    LocalMux I__9666 (
            .O(N__38201),
            .I(N__38198));
    Span4Mux_h I__9665 (
            .O(N__38198),
            .I(N__38195));
    Odrv4 I__9664 (
            .O(N__38195),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_2 ));
    CascadeMux I__9663 (
            .O(N__38192),
            .I(N__38178));
    CascadeMux I__9662 (
            .O(N__38191),
            .I(N__38175));
    CascadeMux I__9661 (
            .O(N__38190),
            .I(N__38169));
    CascadeMux I__9660 (
            .O(N__38189),
            .I(N__38166));
    CascadeMux I__9659 (
            .O(N__38188),
            .I(N__38163));
    CascadeMux I__9658 (
            .O(N__38187),
            .I(N__38160));
    CascadeMux I__9657 (
            .O(N__38186),
            .I(N__38155));
    CascadeMux I__9656 (
            .O(N__38185),
            .I(N__38151));
    CascadeMux I__9655 (
            .O(N__38184),
            .I(N__38148));
    CascadeMux I__9654 (
            .O(N__38183),
            .I(N__38141));
    CascadeMux I__9653 (
            .O(N__38182),
            .I(N__38138));
    CascadeMux I__9652 (
            .O(N__38181),
            .I(N__38133));
    InMux I__9651 (
            .O(N__38178),
            .I(N__38130));
    InMux I__9650 (
            .O(N__38175),
            .I(N__38127));
    CascadeMux I__9649 (
            .O(N__38174),
            .I(N__38124));
    CascadeMux I__9648 (
            .O(N__38173),
            .I(N__38119));
    CascadeMux I__9647 (
            .O(N__38172),
            .I(N__38115));
    InMux I__9646 (
            .O(N__38169),
            .I(N__38112));
    InMux I__9645 (
            .O(N__38166),
            .I(N__38109));
    InMux I__9644 (
            .O(N__38163),
            .I(N__38106));
    InMux I__9643 (
            .O(N__38160),
            .I(N__38103));
    CascadeMux I__9642 (
            .O(N__38159),
            .I(N__38100));
    CascadeMux I__9641 (
            .O(N__38158),
            .I(N__38095));
    InMux I__9640 (
            .O(N__38155),
            .I(N__38092));
    InMux I__9639 (
            .O(N__38154),
            .I(N__38089));
    InMux I__9638 (
            .O(N__38151),
            .I(N__38086));
    InMux I__9637 (
            .O(N__38148),
            .I(N__38083));
    InMux I__9636 (
            .O(N__38147),
            .I(N__38080));
    CascadeMux I__9635 (
            .O(N__38146),
            .I(N__38075));
    CascadeMux I__9634 (
            .O(N__38145),
            .I(N__38072));
    InMux I__9633 (
            .O(N__38144),
            .I(N__38068));
    InMux I__9632 (
            .O(N__38141),
            .I(N__38064));
    InMux I__9631 (
            .O(N__38138),
            .I(N__38061));
    InMux I__9630 (
            .O(N__38137),
            .I(N__38058));
    InMux I__9629 (
            .O(N__38136),
            .I(N__38055));
    InMux I__9628 (
            .O(N__38133),
            .I(N__38052));
    LocalMux I__9627 (
            .O(N__38130),
            .I(N__38047));
    LocalMux I__9626 (
            .O(N__38127),
            .I(N__38047));
    InMux I__9625 (
            .O(N__38124),
            .I(N__38044));
    InMux I__9624 (
            .O(N__38123),
            .I(N__38041));
    InMux I__9623 (
            .O(N__38122),
            .I(N__38038));
    InMux I__9622 (
            .O(N__38119),
            .I(N__38035));
    InMux I__9621 (
            .O(N__38118),
            .I(N__38032));
    InMux I__9620 (
            .O(N__38115),
            .I(N__38029));
    LocalMux I__9619 (
            .O(N__38112),
            .I(N__38026));
    LocalMux I__9618 (
            .O(N__38109),
            .I(N__38019));
    LocalMux I__9617 (
            .O(N__38106),
            .I(N__38019));
    LocalMux I__9616 (
            .O(N__38103),
            .I(N__38019));
    InMux I__9615 (
            .O(N__38100),
            .I(N__38016));
    InMux I__9614 (
            .O(N__38099),
            .I(N__38013));
    InMux I__9613 (
            .O(N__38098),
            .I(N__38010));
    InMux I__9612 (
            .O(N__38095),
            .I(N__38007));
    LocalMux I__9611 (
            .O(N__38092),
            .I(N__38004));
    LocalMux I__9610 (
            .O(N__38089),
            .I(N__37995));
    LocalMux I__9609 (
            .O(N__38086),
            .I(N__37995));
    LocalMux I__9608 (
            .O(N__38083),
            .I(N__37995));
    LocalMux I__9607 (
            .O(N__38080),
            .I(N__37995));
    InMux I__9606 (
            .O(N__38079),
            .I(N__37992));
    InMux I__9605 (
            .O(N__38078),
            .I(N__37989));
    InMux I__9604 (
            .O(N__38075),
            .I(N__37986));
    InMux I__9603 (
            .O(N__38072),
            .I(N__37983));
    InMux I__9602 (
            .O(N__38071),
            .I(N__37980));
    LocalMux I__9601 (
            .O(N__38068),
            .I(N__37977));
    InMux I__9600 (
            .O(N__38067),
            .I(N__37974));
    LocalMux I__9599 (
            .O(N__38064),
            .I(N__37969));
    LocalMux I__9598 (
            .O(N__38061),
            .I(N__37969));
    LocalMux I__9597 (
            .O(N__38058),
            .I(N__37960));
    LocalMux I__9596 (
            .O(N__38055),
            .I(N__37960));
    LocalMux I__9595 (
            .O(N__38052),
            .I(N__37960));
    Span4Mux_v I__9594 (
            .O(N__38047),
            .I(N__37960));
    LocalMux I__9593 (
            .O(N__38044),
            .I(N__37957));
    LocalMux I__9592 (
            .O(N__38041),
            .I(N__37954));
    LocalMux I__9591 (
            .O(N__38038),
            .I(N__37951));
    LocalMux I__9590 (
            .O(N__38035),
            .I(N__37948));
    LocalMux I__9589 (
            .O(N__38032),
            .I(N__37939));
    LocalMux I__9588 (
            .O(N__38029),
            .I(N__37939));
    Span4Mux_s3_h I__9587 (
            .O(N__38026),
            .I(N__37939));
    Span4Mux_v I__9586 (
            .O(N__38019),
            .I(N__37939));
    LocalMux I__9585 (
            .O(N__38016),
            .I(N__37936));
    LocalMux I__9584 (
            .O(N__38013),
            .I(N__37929));
    LocalMux I__9583 (
            .O(N__38010),
            .I(N__37929));
    LocalMux I__9582 (
            .O(N__38007),
            .I(N__37929));
    Span4Mux_v I__9581 (
            .O(N__38004),
            .I(N__37926));
    Span4Mux_v I__9580 (
            .O(N__37995),
            .I(N__37923));
    LocalMux I__9579 (
            .O(N__37992),
            .I(N__37910));
    LocalMux I__9578 (
            .O(N__37989),
            .I(N__37910));
    LocalMux I__9577 (
            .O(N__37986),
            .I(N__37910));
    LocalMux I__9576 (
            .O(N__37983),
            .I(N__37910));
    LocalMux I__9575 (
            .O(N__37980),
            .I(N__37910));
    Span4Mux_s2_v I__9574 (
            .O(N__37977),
            .I(N__37910));
    LocalMux I__9573 (
            .O(N__37974),
            .I(N__37903));
    Span4Mux_v I__9572 (
            .O(N__37969),
            .I(N__37903));
    Span4Mux_v I__9571 (
            .O(N__37960),
            .I(N__37903));
    Span4Mux_s3_h I__9570 (
            .O(N__37957),
            .I(N__37900));
    Span4Mux_v I__9569 (
            .O(N__37954),
            .I(N__37890));
    Span4Mux_s3_h I__9568 (
            .O(N__37951),
            .I(N__37890));
    Span4Mux_v I__9567 (
            .O(N__37948),
            .I(N__37890));
    Span4Mux_v I__9566 (
            .O(N__37939),
            .I(N__37890));
    Span4Mux_v I__9565 (
            .O(N__37936),
            .I(N__37881));
    Span4Mux_v I__9564 (
            .O(N__37929),
            .I(N__37881));
    Span4Mux_h I__9563 (
            .O(N__37926),
            .I(N__37881));
    Span4Mux_h I__9562 (
            .O(N__37923),
            .I(N__37881));
    Span4Mux_v I__9561 (
            .O(N__37910),
            .I(N__37874));
    Span4Mux_h I__9560 (
            .O(N__37903),
            .I(N__37874));
    Span4Mux_v I__9559 (
            .O(N__37900),
            .I(N__37874));
    InMux I__9558 (
            .O(N__37899),
            .I(N__37871));
    Odrv4 I__9557 (
            .O(N__37890),
            .I(\processor_zipi8.arith_logical_result_3 ));
    Odrv4 I__9556 (
            .O(N__37881),
            .I(\processor_zipi8.arith_logical_result_3 ));
    Odrv4 I__9555 (
            .O(N__37874),
            .I(\processor_zipi8.arith_logical_result_3 ));
    LocalMux I__9554 (
            .O(N__37871),
            .I(\processor_zipi8.arith_logical_result_3 ));
    CascadeMux I__9553 (
            .O(N__37862),
            .I(N__37859));
    InMux I__9552 (
            .O(N__37859),
            .I(N__37854));
    CascadeMux I__9551 (
            .O(N__37858),
            .I(N__37850));
    CascadeMux I__9550 (
            .O(N__37857),
            .I(N__37847));
    LocalMux I__9549 (
            .O(N__37854),
            .I(N__37844));
    CascadeMux I__9548 (
            .O(N__37853),
            .I(N__37841));
    InMux I__9547 (
            .O(N__37850),
            .I(N__37837));
    InMux I__9546 (
            .O(N__37847),
            .I(N__37832));
    Span4Mux_v I__9545 (
            .O(N__37844),
            .I(N__37829));
    InMux I__9544 (
            .O(N__37841),
            .I(N__37826));
    CascadeMux I__9543 (
            .O(N__37840),
            .I(N__37820));
    LocalMux I__9542 (
            .O(N__37837),
            .I(N__37817));
    InMux I__9541 (
            .O(N__37836),
            .I(N__37814));
    CascadeMux I__9540 (
            .O(N__37835),
            .I(N__37811));
    LocalMux I__9539 (
            .O(N__37832),
            .I(N__37807));
    Span4Mux_h I__9538 (
            .O(N__37829),
            .I(N__37802));
    LocalMux I__9537 (
            .O(N__37826),
            .I(N__37802));
    InMux I__9536 (
            .O(N__37825),
            .I(N__37798));
    CascadeMux I__9535 (
            .O(N__37824),
            .I(N__37794));
    InMux I__9534 (
            .O(N__37823),
            .I(N__37790));
    InMux I__9533 (
            .O(N__37820),
            .I(N__37787));
    Span4Mux_s0_h I__9532 (
            .O(N__37817),
            .I(N__37782));
    LocalMux I__9531 (
            .O(N__37814),
            .I(N__37782));
    InMux I__9530 (
            .O(N__37811),
            .I(N__37779));
    InMux I__9529 (
            .O(N__37810),
            .I(N__37775));
    Span4Mux_h I__9528 (
            .O(N__37807),
            .I(N__37769));
    Span4Mux_v I__9527 (
            .O(N__37802),
            .I(N__37769));
    InMux I__9526 (
            .O(N__37801),
            .I(N__37766));
    LocalMux I__9525 (
            .O(N__37798),
            .I(N__37763));
    InMux I__9524 (
            .O(N__37797),
            .I(N__37760));
    InMux I__9523 (
            .O(N__37794),
            .I(N__37757));
    InMux I__9522 (
            .O(N__37793),
            .I(N__37750));
    LocalMux I__9521 (
            .O(N__37790),
            .I(N__37741));
    LocalMux I__9520 (
            .O(N__37787),
            .I(N__37741));
    Span4Mux_v I__9519 (
            .O(N__37782),
            .I(N__37741));
    LocalMux I__9518 (
            .O(N__37779),
            .I(N__37741));
    InMux I__9517 (
            .O(N__37778),
            .I(N__37738));
    LocalMux I__9516 (
            .O(N__37775),
            .I(N__37735));
    InMux I__9515 (
            .O(N__37774),
            .I(N__37732));
    Span4Mux_v I__9514 (
            .O(N__37769),
            .I(N__37727));
    LocalMux I__9513 (
            .O(N__37766),
            .I(N__37727));
    Span4Mux_v I__9512 (
            .O(N__37763),
            .I(N__37722));
    LocalMux I__9511 (
            .O(N__37760),
            .I(N__37722));
    LocalMux I__9510 (
            .O(N__37757),
            .I(N__37719));
    InMux I__9509 (
            .O(N__37756),
            .I(N__37716));
    InMux I__9508 (
            .O(N__37755),
            .I(N__37713));
    InMux I__9507 (
            .O(N__37754),
            .I(N__37710));
    InMux I__9506 (
            .O(N__37753),
            .I(N__37707));
    LocalMux I__9505 (
            .O(N__37750),
            .I(N__37698));
    Span4Mux_v I__9504 (
            .O(N__37741),
            .I(N__37693));
    LocalMux I__9503 (
            .O(N__37738),
            .I(N__37693));
    Span4Mux_v I__9502 (
            .O(N__37735),
            .I(N__37690));
    LocalMux I__9501 (
            .O(N__37732),
            .I(N__37685));
    Span4Mux_v I__9500 (
            .O(N__37727),
            .I(N__37685));
    Span4Mux_v I__9499 (
            .O(N__37722),
            .I(N__37680));
    Span4Mux_v I__9498 (
            .O(N__37719),
            .I(N__37680));
    LocalMux I__9497 (
            .O(N__37716),
            .I(N__37677));
    LocalMux I__9496 (
            .O(N__37713),
            .I(N__37674));
    LocalMux I__9495 (
            .O(N__37710),
            .I(N__37669));
    LocalMux I__9494 (
            .O(N__37707),
            .I(N__37669));
    CascadeMux I__9493 (
            .O(N__37706),
            .I(N__37665));
    InMux I__9492 (
            .O(N__37705),
            .I(N__37662));
    CascadeMux I__9491 (
            .O(N__37704),
            .I(N__37658));
    InMux I__9490 (
            .O(N__37703),
            .I(N__37655));
    InMux I__9489 (
            .O(N__37702),
            .I(N__37651));
    InMux I__9488 (
            .O(N__37701),
            .I(N__37648));
    Span4Mux_v I__9487 (
            .O(N__37698),
            .I(N__37641));
    Span4Mux_v I__9486 (
            .O(N__37693),
            .I(N__37641));
    Span4Mux_s0_h I__9485 (
            .O(N__37690),
            .I(N__37641));
    Span4Mux_h I__9484 (
            .O(N__37685),
            .I(N__37630));
    Span4Mux_h I__9483 (
            .O(N__37680),
            .I(N__37630));
    Span4Mux_s2_h I__9482 (
            .O(N__37677),
            .I(N__37630));
    Span4Mux_v I__9481 (
            .O(N__37674),
            .I(N__37630));
    Span4Mux_v I__9480 (
            .O(N__37669),
            .I(N__37630));
    CascadeMux I__9479 (
            .O(N__37668),
            .I(N__37624));
    InMux I__9478 (
            .O(N__37665),
            .I(N__37621));
    LocalMux I__9477 (
            .O(N__37662),
            .I(N__37618));
    InMux I__9476 (
            .O(N__37661),
            .I(N__37615));
    InMux I__9475 (
            .O(N__37658),
            .I(N__37612));
    LocalMux I__9474 (
            .O(N__37655),
            .I(N__37609));
    InMux I__9473 (
            .O(N__37654),
            .I(N__37606));
    LocalMux I__9472 (
            .O(N__37651),
            .I(N__37603));
    LocalMux I__9471 (
            .O(N__37648),
            .I(N__37600));
    Sp12to4 I__9470 (
            .O(N__37641),
            .I(N__37595));
    Sp12to4 I__9469 (
            .O(N__37630),
            .I(N__37595));
    InMux I__9468 (
            .O(N__37629),
            .I(N__37592));
    InMux I__9467 (
            .O(N__37628),
            .I(N__37589));
    InMux I__9466 (
            .O(N__37627),
            .I(N__37586));
    InMux I__9465 (
            .O(N__37624),
            .I(N__37583));
    LocalMux I__9464 (
            .O(N__37621),
            .I(N__37580));
    Span4Mux_s2_v I__9463 (
            .O(N__37618),
            .I(N__37577));
    LocalMux I__9462 (
            .O(N__37615),
            .I(N__37570));
    LocalMux I__9461 (
            .O(N__37612),
            .I(N__37570));
    Span4Mux_v I__9460 (
            .O(N__37609),
            .I(N__37570));
    LocalMux I__9459 (
            .O(N__37606),
            .I(N__37565));
    Span4Mux_v I__9458 (
            .O(N__37603),
            .I(N__37565));
    Span12Mux_s6_h I__9457 (
            .O(N__37600),
            .I(N__37560));
    Span12Mux_s5_h I__9456 (
            .O(N__37595),
            .I(N__37560));
    LocalMux I__9455 (
            .O(N__37592),
            .I(N__37555));
    LocalMux I__9454 (
            .O(N__37589),
            .I(N__37555));
    LocalMux I__9453 (
            .O(N__37586),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    LocalMux I__9452 (
            .O(N__37583),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    Odrv4 I__9451 (
            .O(N__37580),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    Odrv4 I__9450 (
            .O(N__37577),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    Odrv4 I__9449 (
            .O(N__37570),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    Odrv4 I__9448 (
            .O(N__37565),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    Odrv12 I__9447 (
            .O(N__37560),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    Odrv12 I__9446 (
            .O(N__37555),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ));
    InMux I__9445 (
            .O(N__37538),
            .I(N__37535));
    LocalMux I__9444 (
            .O(N__37535),
            .I(N__37531));
    InMux I__9443 (
            .O(N__37534),
            .I(N__37528));
    Span4Mux_v I__9442 (
            .O(N__37531),
            .I(N__37523));
    LocalMux I__9441 (
            .O(N__37528),
            .I(N__37523));
    Span4Mux_s0_h I__9440 (
            .O(N__37523),
            .I(N__37520));
    Odrv4 I__9439 (
            .O(N__37520),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_3 ));
    InMux I__9438 (
            .O(N__37517),
            .I(N__37513));
    InMux I__9437 (
            .O(N__37516),
            .I(N__37510));
    LocalMux I__9436 (
            .O(N__37513),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3 ));
    LocalMux I__9435 (
            .O(N__37510),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3 ));
    InMux I__9434 (
            .O(N__37505),
            .I(N__37491));
    InMux I__9433 (
            .O(N__37504),
            .I(N__37479));
    InMux I__9432 (
            .O(N__37503),
            .I(N__37479));
    InMux I__9431 (
            .O(N__37502),
            .I(N__37470));
    InMux I__9430 (
            .O(N__37501),
            .I(N__37470));
    InMux I__9429 (
            .O(N__37500),
            .I(N__37470));
    InMux I__9428 (
            .O(N__37499),
            .I(N__37462));
    InMux I__9427 (
            .O(N__37498),
            .I(N__37462));
    InMux I__9426 (
            .O(N__37497),
            .I(N__37457));
    InMux I__9425 (
            .O(N__37496),
            .I(N__37457));
    InMux I__9424 (
            .O(N__37495),
            .I(N__37452));
    InMux I__9423 (
            .O(N__37494),
            .I(N__37452));
    LocalMux I__9422 (
            .O(N__37491),
            .I(N__37445));
    InMux I__9421 (
            .O(N__37490),
            .I(N__37442));
    InMux I__9420 (
            .O(N__37489),
            .I(N__37433));
    InMux I__9419 (
            .O(N__37488),
            .I(N__37433));
    InMux I__9418 (
            .O(N__37487),
            .I(N__37420));
    InMux I__9417 (
            .O(N__37486),
            .I(N__37417));
    InMux I__9416 (
            .O(N__37485),
            .I(N__37412));
    InMux I__9415 (
            .O(N__37484),
            .I(N__37412));
    LocalMux I__9414 (
            .O(N__37479),
            .I(N__37406));
    InMux I__9413 (
            .O(N__37478),
            .I(N__37401));
    InMux I__9412 (
            .O(N__37477),
            .I(N__37401));
    LocalMux I__9411 (
            .O(N__37470),
            .I(N__37398));
    InMux I__9410 (
            .O(N__37469),
            .I(N__37391));
    InMux I__9409 (
            .O(N__37468),
            .I(N__37386));
    InMux I__9408 (
            .O(N__37467),
            .I(N__37386));
    LocalMux I__9407 (
            .O(N__37462),
            .I(N__37378));
    LocalMux I__9406 (
            .O(N__37457),
            .I(N__37373));
    LocalMux I__9405 (
            .O(N__37452),
            .I(N__37373));
    InMux I__9404 (
            .O(N__37451),
            .I(N__37369));
    InMux I__9403 (
            .O(N__37450),
            .I(N__37362));
    InMux I__9402 (
            .O(N__37449),
            .I(N__37362));
    InMux I__9401 (
            .O(N__37448),
            .I(N__37362));
    Span4Mux_v I__9400 (
            .O(N__37445),
            .I(N__37357));
    LocalMux I__9399 (
            .O(N__37442),
            .I(N__37357));
    InMux I__9398 (
            .O(N__37441),
            .I(N__37349));
    InMux I__9397 (
            .O(N__37440),
            .I(N__37349));
    InMux I__9396 (
            .O(N__37439),
            .I(N__37346));
    InMux I__9395 (
            .O(N__37438),
            .I(N__37343));
    LocalMux I__9394 (
            .O(N__37433),
            .I(N__37340));
    InMux I__9393 (
            .O(N__37432),
            .I(N__37333));
    InMux I__9392 (
            .O(N__37431),
            .I(N__37333));
    InMux I__9391 (
            .O(N__37430),
            .I(N__37333));
    InMux I__9390 (
            .O(N__37429),
            .I(N__37324));
    InMux I__9389 (
            .O(N__37428),
            .I(N__37317));
    InMux I__9388 (
            .O(N__37427),
            .I(N__37317));
    InMux I__9387 (
            .O(N__37426),
            .I(N__37310));
    InMux I__9386 (
            .O(N__37425),
            .I(N__37310));
    InMux I__9385 (
            .O(N__37424),
            .I(N__37310));
    InMux I__9384 (
            .O(N__37423),
            .I(N__37307));
    LocalMux I__9383 (
            .O(N__37420),
            .I(N__37304));
    LocalMux I__9382 (
            .O(N__37417),
            .I(N__37290));
    LocalMux I__9381 (
            .O(N__37412),
            .I(N__37287));
    InMux I__9380 (
            .O(N__37411),
            .I(N__37281));
    InMux I__9379 (
            .O(N__37410),
            .I(N__37281));
    InMux I__9378 (
            .O(N__37409),
            .I(N__37278));
    Span4Mux_s2_v I__9377 (
            .O(N__37406),
            .I(N__37273));
    LocalMux I__9376 (
            .O(N__37401),
            .I(N__37273));
    Span4Mux_v I__9375 (
            .O(N__37398),
            .I(N__37270));
    InMux I__9374 (
            .O(N__37397),
            .I(N__37265));
    InMux I__9373 (
            .O(N__37396),
            .I(N__37265));
    InMux I__9372 (
            .O(N__37395),
            .I(N__37260));
    InMux I__9371 (
            .O(N__37394),
            .I(N__37260));
    LocalMux I__9370 (
            .O(N__37391),
            .I(N__37255));
    LocalMux I__9369 (
            .O(N__37386),
            .I(N__37255));
    CascadeMux I__9368 (
            .O(N__37385),
            .I(N__37246));
    InMux I__9367 (
            .O(N__37384),
            .I(N__37236));
    InMux I__9366 (
            .O(N__37383),
            .I(N__37236));
    InMux I__9365 (
            .O(N__37382),
            .I(N__37236));
    InMux I__9364 (
            .O(N__37381),
            .I(N__37236));
    Span4Mux_v I__9363 (
            .O(N__37378),
            .I(N__37231));
    Span4Mux_v I__9362 (
            .O(N__37373),
            .I(N__37231));
    InMux I__9361 (
            .O(N__37372),
            .I(N__37228));
    LocalMux I__9360 (
            .O(N__37369),
            .I(N__37221));
    LocalMux I__9359 (
            .O(N__37362),
            .I(N__37221));
    Span4Mux_s3_v I__9358 (
            .O(N__37357),
            .I(N__37221));
    InMux I__9357 (
            .O(N__37356),
            .I(N__37218));
    InMux I__9356 (
            .O(N__37355),
            .I(N__37206));
    InMux I__9355 (
            .O(N__37354),
            .I(N__37206));
    LocalMux I__9354 (
            .O(N__37349),
            .I(N__37203));
    LocalMux I__9353 (
            .O(N__37346),
            .I(N__37194));
    LocalMux I__9352 (
            .O(N__37343),
            .I(N__37194));
    Span4Mux_h I__9351 (
            .O(N__37340),
            .I(N__37194));
    LocalMux I__9350 (
            .O(N__37333),
            .I(N__37194));
    InMux I__9349 (
            .O(N__37332),
            .I(N__37183));
    InMux I__9348 (
            .O(N__37331),
            .I(N__37183));
    InMux I__9347 (
            .O(N__37330),
            .I(N__37183));
    InMux I__9346 (
            .O(N__37329),
            .I(N__37183));
    InMux I__9345 (
            .O(N__37328),
            .I(N__37183));
    InMux I__9344 (
            .O(N__37327),
            .I(N__37180));
    LocalMux I__9343 (
            .O(N__37324),
            .I(N__37177));
    InMux I__9342 (
            .O(N__37323),
            .I(N__37172));
    InMux I__9341 (
            .O(N__37322),
            .I(N__37172));
    LocalMux I__9340 (
            .O(N__37317),
            .I(N__37163));
    LocalMux I__9339 (
            .O(N__37310),
            .I(N__37163));
    LocalMux I__9338 (
            .O(N__37307),
            .I(N__37163));
    Span4Mux_s3_v I__9337 (
            .O(N__37304),
            .I(N__37163));
    InMux I__9336 (
            .O(N__37303),
            .I(N__37154));
    InMux I__9335 (
            .O(N__37302),
            .I(N__37154));
    InMux I__9334 (
            .O(N__37301),
            .I(N__37154));
    InMux I__9333 (
            .O(N__37300),
            .I(N__37154));
    InMux I__9332 (
            .O(N__37299),
            .I(N__37147));
    InMux I__9331 (
            .O(N__37298),
            .I(N__37147));
    InMux I__9330 (
            .O(N__37297),
            .I(N__37147));
    InMux I__9329 (
            .O(N__37296),
            .I(N__37140));
    InMux I__9328 (
            .O(N__37295),
            .I(N__37140));
    InMux I__9327 (
            .O(N__37294),
            .I(N__37140));
    InMux I__9326 (
            .O(N__37293),
            .I(N__37137));
    Span4Mux_v I__9325 (
            .O(N__37290),
            .I(N__37129));
    Span4Mux_h I__9324 (
            .O(N__37287),
            .I(N__37129));
    InMux I__9323 (
            .O(N__37286),
            .I(N__37126));
    LocalMux I__9322 (
            .O(N__37281),
            .I(N__37123));
    LocalMux I__9321 (
            .O(N__37278),
            .I(N__37118));
    Span4Mux_h I__9320 (
            .O(N__37273),
            .I(N__37118));
    IoSpan4Mux I__9319 (
            .O(N__37270),
            .I(N__37113));
    LocalMux I__9318 (
            .O(N__37265),
            .I(N__37113));
    LocalMux I__9317 (
            .O(N__37260),
            .I(N__37108));
    Span4Mux_s3_v I__9316 (
            .O(N__37255),
            .I(N__37108));
    InMux I__9315 (
            .O(N__37254),
            .I(N__37105));
    InMux I__9314 (
            .O(N__37253),
            .I(N__37098));
    InMux I__9313 (
            .O(N__37252),
            .I(N__37098));
    InMux I__9312 (
            .O(N__37251),
            .I(N__37098));
    InMux I__9311 (
            .O(N__37250),
            .I(N__37093));
    InMux I__9310 (
            .O(N__37249),
            .I(N__37093));
    InMux I__9309 (
            .O(N__37246),
            .I(N__37090));
    CascadeMux I__9308 (
            .O(N__37245),
            .I(N__37085));
    LocalMux I__9307 (
            .O(N__37236),
            .I(N__37072));
    Span4Mux_h I__9306 (
            .O(N__37231),
            .I(N__37061));
    LocalMux I__9305 (
            .O(N__37228),
            .I(N__37054));
    Span4Mux_v I__9304 (
            .O(N__37221),
            .I(N__37054));
    LocalMux I__9303 (
            .O(N__37218),
            .I(N__37054));
    InMux I__9302 (
            .O(N__37217),
            .I(N__37049));
    InMux I__9301 (
            .O(N__37216),
            .I(N__37049));
    InMux I__9300 (
            .O(N__37215),
            .I(N__37044));
    InMux I__9299 (
            .O(N__37214),
            .I(N__37044));
    InMux I__9298 (
            .O(N__37213),
            .I(N__37037));
    InMux I__9297 (
            .O(N__37212),
            .I(N__37037));
    InMux I__9296 (
            .O(N__37211),
            .I(N__37037));
    LocalMux I__9295 (
            .O(N__37206),
            .I(N__37034));
    Span4Mux_h I__9294 (
            .O(N__37203),
            .I(N__37029));
    Span4Mux_v I__9293 (
            .O(N__37194),
            .I(N__37029));
    LocalMux I__9292 (
            .O(N__37183),
            .I(N__37012));
    LocalMux I__9291 (
            .O(N__37180),
            .I(N__37012));
    Span4Mux_h I__9290 (
            .O(N__37177),
            .I(N__37012));
    LocalMux I__9289 (
            .O(N__37172),
            .I(N__37012));
    Span4Mux_v I__9288 (
            .O(N__37163),
            .I(N__37012));
    LocalMux I__9287 (
            .O(N__37154),
            .I(N__37012));
    LocalMux I__9286 (
            .O(N__37147),
            .I(N__37012));
    LocalMux I__9285 (
            .O(N__37140),
            .I(N__37012));
    LocalMux I__9284 (
            .O(N__37137),
            .I(N__37009));
    InMux I__9283 (
            .O(N__37136),
            .I(N__37002));
    InMux I__9282 (
            .O(N__37135),
            .I(N__37002));
    InMux I__9281 (
            .O(N__37134),
            .I(N__37002));
    Span4Mux_h I__9280 (
            .O(N__37129),
            .I(N__36991));
    LocalMux I__9279 (
            .O(N__37126),
            .I(N__36991));
    Span4Mux_h I__9278 (
            .O(N__37123),
            .I(N__36991));
    Span4Mux_v I__9277 (
            .O(N__37118),
            .I(N__36991));
    Span4Mux_s2_h I__9276 (
            .O(N__37113),
            .I(N__36991));
    Span4Mux_h I__9275 (
            .O(N__37108),
            .I(N__36986));
    LocalMux I__9274 (
            .O(N__37105),
            .I(N__36986));
    LocalMux I__9273 (
            .O(N__37098),
            .I(N__36983));
    LocalMux I__9272 (
            .O(N__37093),
            .I(N__36980));
    LocalMux I__9271 (
            .O(N__37090),
            .I(N__36977));
    InMux I__9270 (
            .O(N__37089),
            .I(N__36970));
    InMux I__9269 (
            .O(N__37088),
            .I(N__36970));
    InMux I__9268 (
            .O(N__37085),
            .I(N__36970));
    InMux I__9267 (
            .O(N__37084),
            .I(N__36963));
    InMux I__9266 (
            .O(N__37083),
            .I(N__36963));
    InMux I__9265 (
            .O(N__37082),
            .I(N__36963));
    InMux I__9264 (
            .O(N__37081),
            .I(N__36954));
    InMux I__9263 (
            .O(N__37080),
            .I(N__36954));
    InMux I__9262 (
            .O(N__37079),
            .I(N__36954));
    InMux I__9261 (
            .O(N__37078),
            .I(N__36954));
    InMux I__9260 (
            .O(N__37077),
            .I(N__36947));
    InMux I__9259 (
            .O(N__37076),
            .I(N__36947));
    InMux I__9258 (
            .O(N__37075),
            .I(N__36947));
    Span12Mux_s9_h I__9257 (
            .O(N__37072),
            .I(N__36944));
    InMux I__9256 (
            .O(N__37071),
            .I(N__36937));
    InMux I__9255 (
            .O(N__37070),
            .I(N__36937));
    InMux I__9254 (
            .O(N__37069),
            .I(N__36937));
    InMux I__9253 (
            .O(N__37068),
            .I(N__36926));
    InMux I__9252 (
            .O(N__37067),
            .I(N__36926));
    InMux I__9251 (
            .O(N__37066),
            .I(N__36926));
    InMux I__9250 (
            .O(N__37065),
            .I(N__36926));
    InMux I__9249 (
            .O(N__37064),
            .I(N__36926));
    Span4Mux_h I__9248 (
            .O(N__37061),
            .I(N__36919));
    Span4Mux_v I__9247 (
            .O(N__37054),
            .I(N__36919));
    LocalMux I__9246 (
            .O(N__37049),
            .I(N__36919));
    LocalMux I__9245 (
            .O(N__37044),
            .I(N__36908));
    LocalMux I__9244 (
            .O(N__37037),
            .I(N__36908));
    Span4Mux_v I__9243 (
            .O(N__37034),
            .I(N__36908));
    Span4Mux_v I__9242 (
            .O(N__37029),
            .I(N__36908));
    Span4Mux_v I__9241 (
            .O(N__37012),
            .I(N__36908));
    Span4Mux_h I__9240 (
            .O(N__37009),
            .I(N__36901));
    LocalMux I__9239 (
            .O(N__37002),
            .I(N__36901));
    Span4Mux_v I__9238 (
            .O(N__36991),
            .I(N__36901));
    Span4Mux_h I__9237 (
            .O(N__36986),
            .I(N__36890));
    Span4Mux_s2_h I__9236 (
            .O(N__36983),
            .I(N__36890));
    Span4Mux_v I__9235 (
            .O(N__36980),
            .I(N__36890));
    Span4Mux_h I__9234 (
            .O(N__36977),
            .I(N__36890));
    LocalMux I__9233 (
            .O(N__36970),
            .I(N__36890));
    LocalMux I__9232 (
            .O(N__36963),
            .I(N__36885));
    LocalMux I__9231 (
            .O(N__36954),
            .I(N__36885));
    LocalMux I__9230 (
            .O(N__36947),
            .I(instruction_4));
    Odrv12 I__9229 (
            .O(N__36944),
            .I(instruction_4));
    LocalMux I__9228 (
            .O(N__36937),
            .I(instruction_4));
    LocalMux I__9227 (
            .O(N__36926),
            .I(instruction_4));
    Odrv4 I__9226 (
            .O(N__36919),
            .I(instruction_4));
    Odrv4 I__9225 (
            .O(N__36908),
            .I(instruction_4));
    Odrv4 I__9224 (
            .O(N__36901),
            .I(instruction_4));
    Odrv4 I__9223 (
            .O(N__36890),
            .I(instruction_4));
    Odrv12 I__9222 (
            .O(N__36885),
            .I(instruction_4));
    InMux I__9221 (
            .O(N__36866),
            .I(N__36863));
    LocalMux I__9220 (
            .O(N__36863),
            .I(N__36860));
    Span4Mux_v I__9219 (
            .O(N__36860),
            .I(N__36857));
    Odrv4 I__9218 (
            .O(N__36857),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_3 ));
    CascadeMux I__9217 (
            .O(N__36854),
            .I(N__36837));
    CascadeMux I__9216 (
            .O(N__36853),
            .I(N__36826));
    CascadeMux I__9215 (
            .O(N__36852),
            .I(N__36823));
    CascadeMux I__9214 (
            .O(N__36851),
            .I(N__36820));
    InMux I__9213 (
            .O(N__36850),
            .I(N__36815));
    InMux I__9212 (
            .O(N__36849),
            .I(N__36804));
    CascadeMux I__9211 (
            .O(N__36848),
            .I(N__36800));
    InMux I__9210 (
            .O(N__36847),
            .I(N__36775));
    InMux I__9209 (
            .O(N__36846),
            .I(N__36775));
    InMux I__9208 (
            .O(N__36845),
            .I(N__36775));
    InMux I__9207 (
            .O(N__36844),
            .I(N__36775));
    InMux I__9206 (
            .O(N__36843),
            .I(N__36775));
    InMux I__9205 (
            .O(N__36842),
            .I(N__36775));
    InMux I__9204 (
            .O(N__36841),
            .I(N__36775));
    InMux I__9203 (
            .O(N__36840),
            .I(N__36775));
    InMux I__9202 (
            .O(N__36837),
            .I(N__36772));
    InMux I__9201 (
            .O(N__36836),
            .I(N__36761));
    InMux I__9200 (
            .O(N__36835),
            .I(N__36761));
    InMux I__9199 (
            .O(N__36834),
            .I(N__36761));
    InMux I__9198 (
            .O(N__36833),
            .I(N__36761));
    InMux I__9197 (
            .O(N__36832),
            .I(N__36761));
    InMux I__9196 (
            .O(N__36831),
            .I(N__36744));
    InMux I__9195 (
            .O(N__36830),
            .I(N__36744));
    InMux I__9194 (
            .O(N__36829),
            .I(N__36744));
    InMux I__9193 (
            .O(N__36826),
            .I(N__36744));
    InMux I__9192 (
            .O(N__36823),
            .I(N__36744));
    InMux I__9191 (
            .O(N__36820),
            .I(N__36744));
    InMux I__9190 (
            .O(N__36819),
            .I(N__36744));
    InMux I__9189 (
            .O(N__36818),
            .I(N__36744));
    LocalMux I__9188 (
            .O(N__36815),
            .I(N__36733));
    InMux I__9187 (
            .O(N__36814),
            .I(N__36716));
    InMux I__9186 (
            .O(N__36813),
            .I(N__36716));
    InMux I__9185 (
            .O(N__36812),
            .I(N__36716));
    InMux I__9184 (
            .O(N__36811),
            .I(N__36716));
    InMux I__9183 (
            .O(N__36810),
            .I(N__36716));
    InMux I__9182 (
            .O(N__36809),
            .I(N__36716));
    InMux I__9181 (
            .O(N__36808),
            .I(N__36716));
    InMux I__9180 (
            .O(N__36807),
            .I(N__36716));
    LocalMux I__9179 (
            .O(N__36804),
            .I(N__36713));
    CascadeMux I__9178 (
            .O(N__36803),
            .I(N__36702));
    InMux I__9177 (
            .O(N__36800),
            .I(N__36689));
    InMux I__9176 (
            .O(N__36799),
            .I(N__36675));
    InMux I__9175 (
            .O(N__36798),
            .I(N__36675));
    InMux I__9174 (
            .O(N__36797),
            .I(N__36675));
    InMux I__9173 (
            .O(N__36796),
            .I(N__36675));
    InMux I__9172 (
            .O(N__36795),
            .I(N__36675));
    InMux I__9171 (
            .O(N__36794),
            .I(N__36675));
    CascadeMux I__9170 (
            .O(N__36793),
            .I(N__36672));
    CascadeMux I__9169 (
            .O(N__36792),
            .I(N__36669));
    LocalMux I__9168 (
            .O(N__36775),
            .I(N__36652));
    LocalMux I__9167 (
            .O(N__36772),
            .I(N__36645));
    LocalMux I__9166 (
            .O(N__36761),
            .I(N__36645));
    LocalMux I__9165 (
            .O(N__36744),
            .I(N__36645));
    InMux I__9164 (
            .O(N__36743),
            .I(N__36628));
    InMux I__9163 (
            .O(N__36742),
            .I(N__36628));
    InMux I__9162 (
            .O(N__36741),
            .I(N__36628));
    InMux I__9161 (
            .O(N__36740),
            .I(N__36628));
    InMux I__9160 (
            .O(N__36739),
            .I(N__36628));
    InMux I__9159 (
            .O(N__36738),
            .I(N__36628));
    InMux I__9158 (
            .O(N__36737),
            .I(N__36628));
    InMux I__9157 (
            .O(N__36736),
            .I(N__36628));
    Span4Mux_v I__9156 (
            .O(N__36733),
            .I(N__36588));
    LocalMux I__9155 (
            .O(N__36716),
            .I(N__36588));
    Span4Mux_v I__9154 (
            .O(N__36713),
            .I(N__36585));
    InMux I__9153 (
            .O(N__36712),
            .I(N__36568));
    InMux I__9152 (
            .O(N__36711),
            .I(N__36568));
    InMux I__9151 (
            .O(N__36710),
            .I(N__36568));
    InMux I__9150 (
            .O(N__36709),
            .I(N__36568));
    InMux I__9149 (
            .O(N__36708),
            .I(N__36568));
    InMux I__9148 (
            .O(N__36707),
            .I(N__36568));
    InMux I__9147 (
            .O(N__36706),
            .I(N__36568));
    InMux I__9146 (
            .O(N__36705),
            .I(N__36568));
    InMux I__9145 (
            .O(N__36702),
            .I(N__36565));
    CascadeMux I__9144 (
            .O(N__36701),
            .I(N__36562));
    CascadeMux I__9143 (
            .O(N__36700),
            .I(N__36559));
    InMux I__9142 (
            .O(N__36699),
            .I(N__36527));
    InMux I__9141 (
            .O(N__36698),
            .I(N__36527));
    InMux I__9140 (
            .O(N__36697),
            .I(N__36527));
    InMux I__9139 (
            .O(N__36696),
            .I(N__36527));
    InMux I__9138 (
            .O(N__36695),
            .I(N__36527));
    InMux I__9137 (
            .O(N__36694),
            .I(N__36527));
    InMux I__9136 (
            .O(N__36693),
            .I(N__36527));
    InMux I__9135 (
            .O(N__36692),
            .I(N__36527));
    LocalMux I__9134 (
            .O(N__36689),
            .I(N__36519));
    InMux I__9133 (
            .O(N__36688),
            .I(N__36516));
    LocalMux I__9132 (
            .O(N__36675),
            .I(N__36513));
    InMux I__9131 (
            .O(N__36672),
            .I(N__36510));
    InMux I__9130 (
            .O(N__36669),
            .I(N__36507));
    InMux I__9129 (
            .O(N__36668),
            .I(N__36504));
    InMux I__9128 (
            .O(N__36667),
            .I(N__36488));
    InMux I__9127 (
            .O(N__36666),
            .I(N__36488));
    InMux I__9126 (
            .O(N__36665),
            .I(N__36488));
    InMux I__9125 (
            .O(N__36664),
            .I(N__36488));
    InMux I__9124 (
            .O(N__36663),
            .I(N__36488));
    InMux I__9123 (
            .O(N__36662),
            .I(N__36488));
    InMux I__9122 (
            .O(N__36661),
            .I(N__36485));
    InMux I__9121 (
            .O(N__36660),
            .I(N__36477));
    InMux I__9120 (
            .O(N__36659),
            .I(N__36477));
    InMux I__9119 (
            .O(N__36658),
            .I(N__36477));
    InMux I__9118 (
            .O(N__36657),
            .I(N__36470));
    InMux I__9117 (
            .O(N__36656),
            .I(N__36470));
    InMux I__9116 (
            .O(N__36655),
            .I(N__36470));
    Span4Mux_v I__9115 (
            .O(N__36652),
            .I(N__36467));
    Span4Mux_v I__9114 (
            .O(N__36645),
            .I(N__36462));
    LocalMux I__9113 (
            .O(N__36628),
            .I(N__36462));
    CascadeMux I__9112 (
            .O(N__36627),
            .I(N__36459));
    CascadeMux I__9111 (
            .O(N__36626),
            .I(N__36456));
    InMux I__9110 (
            .O(N__36625),
            .I(N__36450));
    InMux I__9109 (
            .O(N__36624),
            .I(N__36450));
    InMux I__9108 (
            .O(N__36623),
            .I(N__36447));
    InMux I__9107 (
            .O(N__36622),
            .I(N__36430));
    InMux I__9106 (
            .O(N__36621),
            .I(N__36430));
    InMux I__9105 (
            .O(N__36620),
            .I(N__36430));
    InMux I__9104 (
            .O(N__36619),
            .I(N__36430));
    InMux I__9103 (
            .O(N__36618),
            .I(N__36430));
    InMux I__9102 (
            .O(N__36617),
            .I(N__36430));
    InMux I__9101 (
            .O(N__36616),
            .I(N__36430));
    InMux I__9100 (
            .O(N__36615),
            .I(N__36430));
    InMux I__9099 (
            .O(N__36614),
            .I(N__36415));
    InMux I__9098 (
            .O(N__36613),
            .I(N__36415));
    InMux I__9097 (
            .O(N__36612),
            .I(N__36415));
    InMux I__9096 (
            .O(N__36611),
            .I(N__36415));
    InMux I__9095 (
            .O(N__36610),
            .I(N__36415));
    InMux I__9094 (
            .O(N__36609),
            .I(N__36415));
    InMux I__9093 (
            .O(N__36608),
            .I(N__36415));
    CascadeMux I__9092 (
            .O(N__36607),
            .I(N__36407));
    CascadeMux I__9091 (
            .O(N__36606),
            .I(N__36400));
    CascadeMux I__9090 (
            .O(N__36605),
            .I(N__36397));
    InMux I__9089 (
            .O(N__36604),
            .I(N__36386));
    InMux I__9088 (
            .O(N__36603),
            .I(N__36386));
    InMux I__9087 (
            .O(N__36602),
            .I(N__36386));
    InMux I__9086 (
            .O(N__36601),
            .I(N__36386));
    InMux I__9085 (
            .O(N__36600),
            .I(N__36386));
    CascadeMux I__9084 (
            .O(N__36599),
            .I(N__36374));
    InMux I__9083 (
            .O(N__36598),
            .I(N__36353));
    InMux I__9082 (
            .O(N__36597),
            .I(N__36353));
    InMux I__9081 (
            .O(N__36596),
            .I(N__36353));
    InMux I__9080 (
            .O(N__36595),
            .I(N__36353));
    InMux I__9079 (
            .O(N__36594),
            .I(N__36353));
    InMux I__9078 (
            .O(N__36593),
            .I(N__36353));
    Span4Mux_h I__9077 (
            .O(N__36588),
            .I(N__36344));
    Span4Mux_h I__9076 (
            .O(N__36585),
            .I(N__36344));
    LocalMux I__9075 (
            .O(N__36568),
            .I(N__36344));
    LocalMux I__9074 (
            .O(N__36565),
            .I(N__36344));
    InMux I__9073 (
            .O(N__36562),
            .I(N__36341));
    InMux I__9072 (
            .O(N__36559),
            .I(N__36338));
    InMux I__9071 (
            .O(N__36558),
            .I(N__36333));
    InMux I__9070 (
            .O(N__36557),
            .I(N__36333));
    InMux I__9069 (
            .O(N__36556),
            .I(N__36316));
    InMux I__9068 (
            .O(N__36555),
            .I(N__36316));
    InMux I__9067 (
            .O(N__36554),
            .I(N__36316));
    InMux I__9066 (
            .O(N__36553),
            .I(N__36316));
    InMux I__9065 (
            .O(N__36552),
            .I(N__36316));
    InMux I__9064 (
            .O(N__36551),
            .I(N__36316));
    InMux I__9063 (
            .O(N__36550),
            .I(N__36316));
    InMux I__9062 (
            .O(N__36549),
            .I(N__36316));
    InMux I__9061 (
            .O(N__36548),
            .I(N__36298));
    InMux I__9060 (
            .O(N__36547),
            .I(N__36298));
    InMux I__9059 (
            .O(N__36546),
            .I(N__36298));
    InMux I__9058 (
            .O(N__36545),
            .I(N__36298));
    InMux I__9057 (
            .O(N__36544),
            .I(N__36298));
    LocalMux I__9056 (
            .O(N__36527),
            .I(N__36295));
    InMux I__9055 (
            .O(N__36526),
            .I(N__36288));
    InMux I__9054 (
            .O(N__36525),
            .I(N__36288));
    InMux I__9053 (
            .O(N__36524),
            .I(N__36288));
    CascadeMux I__9052 (
            .O(N__36523),
            .I(N__36285));
    CascadeMux I__9051 (
            .O(N__36522),
            .I(N__36276));
    Span4Mux_v I__9050 (
            .O(N__36519),
            .I(N__36263));
    LocalMux I__9049 (
            .O(N__36516),
            .I(N__36263));
    Span4Mux_v I__9048 (
            .O(N__36513),
            .I(N__36263));
    LocalMux I__9047 (
            .O(N__36510),
            .I(N__36263));
    LocalMux I__9046 (
            .O(N__36507),
            .I(N__36263));
    LocalMux I__9045 (
            .O(N__36504),
            .I(N__36263));
    InMux I__9044 (
            .O(N__36503),
            .I(N__36258));
    InMux I__9043 (
            .O(N__36502),
            .I(N__36258));
    InMux I__9042 (
            .O(N__36501),
            .I(N__36255));
    LocalMux I__9041 (
            .O(N__36488),
            .I(N__36252));
    LocalMux I__9040 (
            .O(N__36485),
            .I(N__36249));
    InMux I__9039 (
            .O(N__36484),
            .I(N__36246));
    LocalMux I__9038 (
            .O(N__36477),
            .I(N__36237));
    LocalMux I__9037 (
            .O(N__36470),
            .I(N__36237));
    Span4Mux_s0_h I__9036 (
            .O(N__36467),
            .I(N__36237));
    Span4Mux_v I__9035 (
            .O(N__36462),
            .I(N__36237));
    InMux I__9034 (
            .O(N__36459),
            .I(N__36234));
    InMux I__9033 (
            .O(N__36456),
            .I(N__36231));
    InMux I__9032 (
            .O(N__36455),
            .I(N__36228));
    LocalMux I__9031 (
            .O(N__36450),
            .I(N__36223));
    LocalMux I__9030 (
            .O(N__36447),
            .I(N__36223));
    LocalMux I__9029 (
            .O(N__36430),
            .I(N__36218));
    LocalMux I__9028 (
            .O(N__36415),
            .I(N__36218));
    InMux I__9027 (
            .O(N__36414),
            .I(N__36207));
    InMux I__9026 (
            .O(N__36413),
            .I(N__36207));
    InMux I__9025 (
            .O(N__36412),
            .I(N__36207));
    InMux I__9024 (
            .O(N__36411),
            .I(N__36207));
    InMux I__9023 (
            .O(N__36410),
            .I(N__36207));
    InMux I__9022 (
            .O(N__36407),
            .I(N__36204));
    InMux I__9021 (
            .O(N__36406),
            .I(N__36168));
    InMux I__9020 (
            .O(N__36405),
            .I(N__36168));
    InMux I__9019 (
            .O(N__36404),
            .I(N__36168));
    InMux I__9018 (
            .O(N__36403),
            .I(N__36168));
    InMux I__9017 (
            .O(N__36400),
            .I(N__36168));
    InMux I__9016 (
            .O(N__36397),
            .I(N__36168));
    LocalMux I__9015 (
            .O(N__36386),
            .I(N__36165));
    InMux I__9014 (
            .O(N__36385),
            .I(N__36148));
    InMux I__9013 (
            .O(N__36384),
            .I(N__36148));
    InMux I__9012 (
            .O(N__36383),
            .I(N__36148));
    InMux I__9011 (
            .O(N__36382),
            .I(N__36148));
    InMux I__9010 (
            .O(N__36381),
            .I(N__36148));
    InMux I__9009 (
            .O(N__36380),
            .I(N__36148));
    InMux I__9008 (
            .O(N__36379),
            .I(N__36148));
    InMux I__9007 (
            .O(N__36378),
            .I(N__36148));
    InMux I__9006 (
            .O(N__36377),
            .I(N__36145));
    InMux I__9005 (
            .O(N__36374),
            .I(N__36134));
    InMux I__9004 (
            .O(N__36373),
            .I(N__36117));
    InMux I__9003 (
            .O(N__36372),
            .I(N__36117));
    InMux I__9002 (
            .O(N__36371),
            .I(N__36117));
    InMux I__9001 (
            .O(N__36370),
            .I(N__36117));
    InMux I__9000 (
            .O(N__36369),
            .I(N__36117));
    InMux I__8999 (
            .O(N__36368),
            .I(N__36117));
    InMux I__8998 (
            .O(N__36367),
            .I(N__36117));
    InMux I__8997 (
            .O(N__36366),
            .I(N__36117));
    LocalMux I__8996 (
            .O(N__36353),
            .I(N__36112));
    Span4Mux_v I__8995 (
            .O(N__36344),
            .I(N__36112));
    LocalMux I__8994 (
            .O(N__36341),
            .I(N__36103));
    LocalMux I__8993 (
            .O(N__36338),
            .I(N__36103));
    LocalMux I__8992 (
            .O(N__36333),
            .I(N__36103));
    LocalMux I__8991 (
            .O(N__36316),
            .I(N__36103));
    InMux I__8990 (
            .O(N__36315),
            .I(N__36095));
    InMux I__8989 (
            .O(N__36314),
            .I(N__36082));
    InMux I__8988 (
            .O(N__36313),
            .I(N__36082));
    InMux I__8987 (
            .O(N__36312),
            .I(N__36082));
    InMux I__8986 (
            .O(N__36311),
            .I(N__36082));
    InMux I__8985 (
            .O(N__36310),
            .I(N__36082));
    InMux I__8984 (
            .O(N__36309),
            .I(N__36082));
    LocalMux I__8983 (
            .O(N__36298),
            .I(N__36079));
    Span4Mux_v I__8982 (
            .O(N__36295),
            .I(N__36074));
    LocalMux I__8981 (
            .O(N__36288),
            .I(N__36074));
    InMux I__8980 (
            .O(N__36285),
            .I(N__36071));
    InMux I__8979 (
            .O(N__36284),
            .I(N__36058));
    InMux I__8978 (
            .O(N__36283),
            .I(N__36058));
    InMux I__8977 (
            .O(N__36282),
            .I(N__36058));
    InMux I__8976 (
            .O(N__36281),
            .I(N__36058));
    InMux I__8975 (
            .O(N__36280),
            .I(N__36058));
    InMux I__8974 (
            .O(N__36279),
            .I(N__36058));
    InMux I__8973 (
            .O(N__36276),
            .I(N__36055));
    Span4Mux_h I__8972 (
            .O(N__36263),
            .I(N__36052));
    LocalMux I__8971 (
            .O(N__36258),
            .I(N__36035));
    LocalMux I__8970 (
            .O(N__36255),
            .I(N__36035));
    Span4Mux_v I__8969 (
            .O(N__36252),
            .I(N__36035));
    Span4Mux_s3_h I__8968 (
            .O(N__36249),
            .I(N__36035));
    LocalMux I__8967 (
            .O(N__36246),
            .I(N__36035));
    Span4Mux_h I__8966 (
            .O(N__36237),
            .I(N__36035));
    LocalMux I__8965 (
            .O(N__36234),
            .I(N__36035));
    LocalMux I__8964 (
            .O(N__36231),
            .I(N__36029));
    LocalMux I__8963 (
            .O(N__36228),
            .I(N__36029));
    Span4Mux_s3_v I__8962 (
            .O(N__36223),
            .I(N__36024));
    Span4Mux_h I__8961 (
            .O(N__36218),
            .I(N__36024));
    LocalMux I__8960 (
            .O(N__36207),
            .I(N__36019));
    LocalMux I__8959 (
            .O(N__36204),
            .I(N__36019));
    InMux I__8958 (
            .O(N__36203),
            .I(N__36002));
    InMux I__8957 (
            .O(N__36202),
            .I(N__36002));
    InMux I__8956 (
            .O(N__36201),
            .I(N__36002));
    InMux I__8955 (
            .O(N__36200),
            .I(N__36002));
    InMux I__8954 (
            .O(N__36199),
            .I(N__36002));
    InMux I__8953 (
            .O(N__36198),
            .I(N__36002));
    InMux I__8952 (
            .O(N__36197),
            .I(N__36002));
    InMux I__8951 (
            .O(N__36196),
            .I(N__36002));
    CascadeMux I__8950 (
            .O(N__36195),
            .I(N__35999));
    CascadeMux I__8949 (
            .O(N__36194),
            .I(N__35996));
    InMux I__8948 (
            .O(N__36193),
            .I(N__35952));
    InMux I__8947 (
            .O(N__36192),
            .I(N__35952));
    InMux I__8946 (
            .O(N__36191),
            .I(N__35952));
    InMux I__8945 (
            .O(N__36190),
            .I(N__35952));
    InMux I__8944 (
            .O(N__36189),
            .I(N__35952));
    InMux I__8943 (
            .O(N__36188),
            .I(N__35952));
    InMux I__8942 (
            .O(N__36187),
            .I(N__35952));
    InMux I__8941 (
            .O(N__36186),
            .I(N__35952));
    InMux I__8940 (
            .O(N__36185),
            .I(N__35941));
    InMux I__8939 (
            .O(N__36184),
            .I(N__35941));
    InMux I__8938 (
            .O(N__36183),
            .I(N__35941));
    InMux I__8937 (
            .O(N__36182),
            .I(N__35941));
    InMux I__8936 (
            .O(N__36181),
            .I(N__35941));
    LocalMux I__8935 (
            .O(N__36168),
            .I(N__35934));
    Span4Mux_v I__8934 (
            .O(N__36165),
            .I(N__35934));
    LocalMux I__8933 (
            .O(N__36148),
            .I(N__35934));
    LocalMux I__8932 (
            .O(N__36145),
            .I(N__35931));
    InMux I__8931 (
            .O(N__36144),
            .I(N__35926));
    InMux I__8930 (
            .O(N__36143),
            .I(N__35926));
    InMux I__8929 (
            .O(N__36142),
            .I(N__35913));
    InMux I__8928 (
            .O(N__36141),
            .I(N__35913));
    InMux I__8927 (
            .O(N__36140),
            .I(N__35913));
    InMux I__8926 (
            .O(N__36139),
            .I(N__35913));
    InMux I__8925 (
            .O(N__36138),
            .I(N__35913));
    InMux I__8924 (
            .O(N__36137),
            .I(N__35913));
    LocalMux I__8923 (
            .O(N__36134),
            .I(N__35910));
    LocalMux I__8922 (
            .O(N__36117),
            .I(N__35907));
    Span4Mux_h I__8921 (
            .O(N__36112),
            .I(N__35902));
    Span4Mux_v I__8920 (
            .O(N__36103),
            .I(N__35902));
    InMux I__8919 (
            .O(N__36102),
            .I(N__35899));
    InMux I__8918 (
            .O(N__36101),
            .I(N__35896));
    CascadeMux I__8917 (
            .O(N__36100),
            .I(N__35893));
    CascadeMux I__8916 (
            .O(N__36099),
            .I(N__35890));
    CascadeMux I__8915 (
            .O(N__36098),
            .I(N__35887));
    LocalMux I__8914 (
            .O(N__36095),
            .I(N__35871));
    LocalMux I__8913 (
            .O(N__36082),
            .I(N__35871));
    Span4Mux_s3_h I__8912 (
            .O(N__36079),
            .I(N__35862));
    Span4Mux_h I__8911 (
            .O(N__36074),
            .I(N__35862));
    LocalMux I__8910 (
            .O(N__36071),
            .I(N__35862));
    LocalMux I__8909 (
            .O(N__36058),
            .I(N__35862));
    LocalMux I__8908 (
            .O(N__36055),
            .I(N__35854));
    Span4Mux_h I__8907 (
            .O(N__36052),
            .I(N__35854));
    InMux I__8906 (
            .O(N__36051),
            .I(N__35849));
    InMux I__8905 (
            .O(N__36050),
            .I(N__35849));
    Span4Mux_h I__8904 (
            .O(N__36035),
            .I(N__35840));
    InMux I__8903 (
            .O(N__36034),
            .I(N__35837));
    Span4Mux_s3_v I__8902 (
            .O(N__36029),
            .I(N__35832));
    Span4Mux_h I__8901 (
            .O(N__36024),
            .I(N__35832));
    Span4Mux_h I__8900 (
            .O(N__36019),
            .I(N__35827));
    LocalMux I__8899 (
            .O(N__36002),
            .I(N__35827));
    InMux I__8898 (
            .O(N__35999),
            .I(N__35822));
    InMux I__8897 (
            .O(N__35996),
            .I(N__35822));
    InMux I__8896 (
            .O(N__35995),
            .I(N__35809));
    InMux I__8895 (
            .O(N__35994),
            .I(N__35809));
    InMux I__8894 (
            .O(N__35993),
            .I(N__35809));
    InMux I__8893 (
            .O(N__35992),
            .I(N__35809));
    InMux I__8892 (
            .O(N__35991),
            .I(N__35809));
    InMux I__8891 (
            .O(N__35990),
            .I(N__35809));
    InMux I__8890 (
            .O(N__35989),
            .I(N__35798));
    InMux I__8889 (
            .O(N__35988),
            .I(N__35798));
    InMux I__8888 (
            .O(N__35987),
            .I(N__35798));
    InMux I__8887 (
            .O(N__35986),
            .I(N__35798));
    InMux I__8886 (
            .O(N__35985),
            .I(N__35798));
    InMux I__8885 (
            .O(N__35984),
            .I(N__35791));
    InMux I__8884 (
            .O(N__35983),
            .I(N__35791));
    InMux I__8883 (
            .O(N__35982),
            .I(N__35791));
    InMux I__8882 (
            .O(N__35981),
            .I(N__35778));
    InMux I__8881 (
            .O(N__35980),
            .I(N__35778));
    InMux I__8880 (
            .O(N__35979),
            .I(N__35778));
    InMux I__8879 (
            .O(N__35978),
            .I(N__35778));
    InMux I__8878 (
            .O(N__35977),
            .I(N__35778));
    InMux I__8877 (
            .O(N__35976),
            .I(N__35778));
    InMux I__8876 (
            .O(N__35975),
            .I(N__35763));
    InMux I__8875 (
            .O(N__35974),
            .I(N__35763));
    InMux I__8874 (
            .O(N__35973),
            .I(N__35763));
    InMux I__8873 (
            .O(N__35972),
            .I(N__35763));
    InMux I__8872 (
            .O(N__35971),
            .I(N__35763));
    InMux I__8871 (
            .O(N__35970),
            .I(N__35763));
    InMux I__8870 (
            .O(N__35969),
            .I(N__35763));
    LocalMux I__8869 (
            .O(N__35952),
            .I(N__35758));
    LocalMux I__8868 (
            .O(N__35941),
            .I(N__35758));
    Span4Mux_h I__8867 (
            .O(N__35934),
            .I(N__35755));
    Span4Mux_v I__8866 (
            .O(N__35931),
            .I(N__35750));
    LocalMux I__8865 (
            .O(N__35926),
            .I(N__35750));
    LocalMux I__8864 (
            .O(N__35913),
            .I(N__35747));
    Span4Mux_v I__8863 (
            .O(N__35910),
            .I(N__35742));
    Span4Mux_v I__8862 (
            .O(N__35907),
            .I(N__35737));
    Span4Mux_v I__8861 (
            .O(N__35902),
            .I(N__35737));
    LocalMux I__8860 (
            .O(N__35899),
            .I(N__35732));
    LocalMux I__8859 (
            .O(N__35896),
            .I(N__35732));
    InMux I__8858 (
            .O(N__35893),
            .I(N__35727));
    InMux I__8857 (
            .O(N__35890),
            .I(N__35724));
    InMux I__8856 (
            .O(N__35887),
            .I(N__35715));
    InMux I__8855 (
            .O(N__35886),
            .I(N__35715));
    InMux I__8854 (
            .O(N__35885),
            .I(N__35715));
    InMux I__8853 (
            .O(N__35884),
            .I(N__35715));
    InMux I__8852 (
            .O(N__35883),
            .I(N__35698));
    InMux I__8851 (
            .O(N__35882),
            .I(N__35698));
    InMux I__8850 (
            .O(N__35881),
            .I(N__35698));
    InMux I__8849 (
            .O(N__35880),
            .I(N__35698));
    InMux I__8848 (
            .O(N__35879),
            .I(N__35698));
    InMux I__8847 (
            .O(N__35878),
            .I(N__35698));
    InMux I__8846 (
            .O(N__35877),
            .I(N__35698));
    InMux I__8845 (
            .O(N__35876),
            .I(N__35698));
    Span4Mux_s2_v I__8844 (
            .O(N__35871),
            .I(N__35693));
    Span4Mux_v I__8843 (
            .O(N__35862),
            .I(N__35693));
    InMux I__8842 (
            .O(N__35861),
            .I(N__35686));
    InMux I__8841 (
            .O(N__35860),
            .I(N__35686));
    InMux I__8840 (
            .O(N__35859),
            .I(N__35686));
    Sp12to4 I__8839 (
            .O(N__35854),
            .I(N__35681));
    LocalMux I__8838 (
            .O(N__35849),
            .I(N__35681));
    InMux I__8837 (
            .O(N__35848),
            .I(N__35668));
    InMux I__8836 (
            .O(N__35847),
            .I(N__35668));
    InMux I__8835 (
            .O(N__35846),
            .I(N__35668));
    InMux I__8834 (
            .O(N__35845),
            .I(N__35668));
    InMux I__8833 (
            .O(N__35844),
            .I(N__35668));
    InMux I__8832 (
            .O(N__35843),
            .I(N__35668));
    Sp12to4 I__8831 (
            .O(N__35840),
            .I(N__35663));
    LocalMux I__8830 (
            .O(N__35837),
            .I(N__35663));
    Span4Mux_v I__8829 (
            .O(N__35832),
            .I(N__35658));
    Span4Mux_s3_h I__8828 (
            .O(N__35827),
            .I(N__35658));
    LocalMux I__8827 (
            .O(N__35822),
            .I(N__35649));
    LocalMux I__8826 (
            .O(N__35809),
            .I(N__35649));
    LocalMux I__8825 (
            .O(N__35798),
            .I(N__35649));
    LocalMux I__8824 (
            .O(N__35791),
            .I(N__35649));
    LocalMux I__8823 (
            .O(N__35778),
            .I(N__35644));
    LocalMux I__8822 (
            .O(N__35763),
            .I(N__35644));
    Span4Mux_h I__8821 (
            .O(N__35758),
            .I(N__35637));
    Span4Mux_v I__8820 (
            .O(N__35755),
            .I(N__35637));
    Span4Mux_v I__8819 (
            .O(N__35750),
            .I(N__35637));
    Span4Mux_h I__8818 (
            .O(N__35747),
            .I(N__35634));
    InMux I__8817 (
            .O(N__35746),
            .I(N__35629));
    InMux I__8816 (
            .O(N__35745),
            .I(N__35629));
    Span4Mux_h I__8815 (
            .O(N__35742),
            .I(N__35622));
    Span4Mux_v I__8814 (
            .O(N__35737),
            .I(N__35622));
    Span4Mux_s2_v I__8813 (
            .O(N__35732),
            .I(N__35622));
    InMux I__8812 (
            .O(N__35731),
            .I(N__35617));
    InMux I__8811 (
            .O(N__35730),
            .I(N__35617));
    LocalMux I__8810 (
            .O(N__35727),
            .I(N__35600));
    LocalMux I__8809 (
            .O(N__35724),
            .I(N__35600));
    LocalMux I__8808 (
            .O(N__35715),
            .I(N__35600));
    LocalMux I__8807 (
            .O(N__35698),
            .I(N__35600));
    Sp12to4 I__8806 (
            .O(N__35693),
            .I(N__35600));
    LocalMux I__8805 (
            .O(N__35686),
            .I(N__35600));
    Span12Mux_v I__8804 (
            .O(N__35681),
            .I(N__35600));
    LocalMux I__8803 (
            .O(N__35668),
            .I(N__35600));
    Span12Mux_s8_v I__8802 (
            .O(N__35663),
            .I(N__35593));
    Sp12to4 I__8801 (
            .O(N__35658),
            .I(N__35593));
    Span12Mux_s8_h I__8800 (
            .O(N__35649),
            .I(N__35593));
    Span4Mux_h I__8799 (
            .O(N__35644),
            .I(N__35588));
    Span4Mux_h I__8798 (
            .O(N__35637),
            .I(N__35588));
    Odrv4 I__8797 (
            .O(N__35634),
            .I(\processor_zipi8.alu_mux_sel_1 ));
    LocalMux I__8796 (
            .O(N__35629),
            .I(\processor_zipi8.alu_mux_sel_1 ));
    Odrv4 I__8795 (
            .O(N__35622),
            .I(\processor_zipi8.alu_mux_sel_1 ));
    LocalMux I__8794 (
            .O(N__35617),
            .I(\processor_zipi8.alu_mux_sel_1 ));
    Odrv12 I__8793 (
            .O(N__35600),
            .I(\processor_zipi8.alu_mux_sel_1 ));
    Odrv12 I__8792 (
            .O(N__35593),
            .I(\processor_zipi8.alu_mux_sel_1 ));
    Odrv4 I__8791 (
            .O(N__35588),
            .I(\processor_zipi8.alu_mux_sel_1 ));
    InMux I__8790 (
            .O(N__35573),
            .I(N__35570));
    LocalMux I__8789 (
            .O(N__35570),
            .I(N__35564));
    CascadeMux I__8788 (
            .O(N__35569),
            .I(N__35561));
    CascadeMux I__8787 (
            .O(N__35568),
            .I(N__35553));
    CascadeMux I__8786 (
            .O(N__35567),
            .I(N__35550));
    Span4Mux_v I__8785 (
            .O(N__35564),
            .I(N__35542));
    InMux I__8784 (
            .O(N__35561),
            .I(N__35539));
    CascadeMux I__8783 (
            .O(N__35560),
            .I(N__35536));
    CascadeMux I__8782 (
            .O(N__35559),
            .I(N__35532));
    CascadeMux I__8781 (
            .O(N__35558),
            .I(N__35527));
    CascadeMux I__8780 (
            .O(N__35557),
            .I(N__35524));
    CascadeMux I__8779 (
            .O(N__35556),
            .I(N__35518));
    InMux I__8778 (
            .O(N__35553),
            .I(N__35515));
    InMux I__8777 (
            .O(N__35550),
            .I(N__35512));
    InMux I__8776 (
            .O(N__35549),
            .I(N__35508));
    CascadeMux I__8775 (
            .O(N__35548),
            .I(N__35505));
    InMux I__8774 (
            .O(N__35547),
            .I(N__35502));
    InMux I__8773 (
            .O(N__35546),
            .I(N__35499));
    InMux I__8772 (
            .O(N__35545),
            .I(N__35495));
    Span4Mux_s2_h I__8771 (
            .O(N__35542),
            .I(N__35489));
    LocalMux I__8770 (
            .O(N__35539),
            .I(N__35489));
    InMux I__8769 (
            .O(N__35536),
            .I(N__35486));
    CascadeMux I__8768 (
            .O(N__35535),
            .I(N__35482));
    InMux I__8767 (
            .O(N__35532),
            .I(N__35479));
    InMux I__8766 (
            .O(N__35531),
            .I(N__35476));
    InMux I__8765 (
            .O(N__35530),
            .I(N__35473));
    InMux I__8764 (
            .O(N__35527),
            .I(N__35469));
    InMux I__8763 (
            .O(N__35524),
            .I(N__35466));
    InMux I__8762 (
            .O(N__35523),
            .I(N__35463));
    InMux I__8761 (
            .O(N__35522),
            .I(N__35460));
    InMux I__8760 (
            .O(N__35521),
            .I(N__35457));
    InMux I__8759 (
            .O(N__35518),
            .I(N__35454));
    LocalMux I__8758 (
            .O(N__35515),
            .I(N__35449));
    LocalMux I__8757 (
            .O(N__35512),
            .I(N__35449));
    InMux I__8756 (
            .O(N__35511),
            .I(N__35446));
    LocalMux I__8755 (
            .O(N__35508),
            .I(N__35443));
    InMux I__8754 (
            .O(N__35505),
            .I(N__35440));
    LocalMux I__8753 (
            .O(N__35502),
            .I(N__35435));
    LocalMux I__8752 (
            .O(N__35499),
            .I(N__35435));
    InMux I__8751 (
            .O(N__35498),
            .I(N__35432));
    LocalMux I__8750 (
            .O(N__35495),
            .I(N__35429));
    InMux I__8749 (
            .O(N__35494),
            .I(N__35423));
    Span4Mux_v I__8748 (
            .O(N__35489),
            .I(N__35418));
    LocalMux I__8747 (
            .O(N__35486),
            .I(N__35418));
    InMux I__8746 (
            .O(N__35485),
            .I(N__35415));
    InMux I__8745 (
            .O(N__35482),
            .I(N__35410));
    LocalMux I__8744 (
            .O(N__35479),
            .I(N__35405));
    LocalMux I__8743 (
            .O(N__35476),
            .I(N__35405));
    LocalMux I__8742 (
            .O(N__35473),
            .I(N__35402));
    InMux I__8741 (
            .O(N__35472),
            .I(N__35399));
    LocalMux I__8740 (
            .O(N__35469),
            .I(N__35396));
    LocalMux I__8739 (
            .O(N__35466),
            .I(N__35393));
    LocalMux I__8738 (
            .O(N__35463),
            .I(N__35382));
    LocalMux I__8737 (
            .O(N__35460),
            .I(N__35382));
    LocalMux I__8736 (
            .O(N__35457),
            .I(N__35382));
    LocalMux I__8735 (
            .O(N__35454),
            .I(N__35382));
    Span4Mux_s2_v I__8734 (
            .O(N__35449),
            .I(N__35382));
    LocalMux I__8733 (
            .O(N__35446),
            .I(N__35377));
    Span4Mux_v I__8732 (
            .O(N__35443),
            .I(N__35377));
    LocalMux I__8731 (
            .O(N__35440),
            .I(N__35372));
    Span4Mux_v I__8730 (
            .O(N__35435),
            .I(N__35372));
    LocalMux I__8729 (
            .O(N__35432),
            .I(N__35367));
    Span4Mux_s1_h I__8728 (
            .O(N__35429),
            .I(N__35367));
    InMux I__8727 (
            .O(N__35428),
            .I(N__35364));
    InMux I__8726 (
            .O(N__35427),
            .I(N__35360));
    InMux I__8725 (
            .O(N__35426),
            .I(N__35357));
    LocalMux I__8724 (
            .O(N__35423),
            .I(N__35354));
    Span4Mux_v I__8723 (
            .O(N__35418),
            .I(N__35351));
    LocalMux I__8722 (
            .O(N__35415),
            .I(N__35348));
    InMux I__8721 (
            .O(N__35414),
            .I(N__35344));
    CascadeMux I__8720 (
            .O(N__35413),
            .I(N__35341));
    LocalMux I__8719 (
            .O(N__35410),
            .I(N__35333));
    Span4Mux_s1_h I__8718 (
            .O(N__35405),
            .I(N__35333));
    Span4Mux_v I__8717 (
            .O(N__35402),
            .I(N__35333));
    LocalMux I__8716 (
            .O(N__35399),
            .I(N__35328));
    Span4Mux_s1_h I__8715 (
            .O(N__35396),
            .I(N__35328));
    Span4Mux_s3_h I__8714 (
            .O(N__35393),
            .I(N__35319));
    Span4Mux_v I__8713 (
            .O(N__35382),
            .I(N__35319));
    Span4Mux_v I__8712 (
            .O(N__35377),
            .I(N__35319));
    Span4Mux_v I__8711 (
            .O(N__35372),
            .I(N__35319));
    Sp12to4 I__8710 (
            .O(N__35367),
            .I(N__35314));
    LocalMux I__8709 (
            .O(N__35364),
            .I(N__35314));
    InMux I__8708 (
            .O(N__35363),
            .I(N__35311));
    LocalMux I__8707 (
            .O(N__35360),
            .I(N__35306));
    LocalMux I__8706 (
            .O(N__35357),
            .I(N__35306));
    Span4Mux_v I__8705 (
            .O(N__35354),
            .I(N__35303));
    Span4Mux_h I__8704 (
            .O(N__35351),
            .I(N__35298));
    Span4Mux_s1_h I__8703 (
            .O(N__35348),
            .I(N__35298));
    InMux I__8702 (
            .O(N__35347),
            .I(N__35294));
    LocalMux I__8701 (
            .O(N__35344),
            .I(N__35291));
    InMux I__8700 (
            .O(N__35341),
            .I(N__35288));
    InMux I__8699 (
            .O(N__35340),
            .I(N__35285));
    Span4Mux_h I__8698 (
            .O(N__35333),
            .I(N__35280));
    Span4Mux_h I__8697 (
            .O(N__35328),
            .I(N__35280));
    Sp12to4 I__8696 (
            .O(N__35319),
            .I(N__35275));
    Span12Mux_s9_v I__8695 (
            .O(N__35314),
            .I(N__35275));
    LocalMux I__8694 (
            .O(N__35311),
            .I(N__35268));
    Span4Mux_v I__8693 (
            .O(N__35306),
            .I(N__35268));
    Span4Mux_h I__8692 (
            .O(N__35303),
            .I(N__35268));
    Span4Mux_h I__8691 (
            .O(N__35298),
            .I(N__35265));
    InMux I__8690 (
            .O(N__35297),
            .I(N__35262));
    LocalMux I__8689 (
            .O(N__35294),
            .I(N__35255));
    Span12Mux_s6_h I__8688 (
            .O(N__35291),
            .I(N__35255));
    LocalMux I__8687 (
            .O(N__35288),
            .I(N__35255));
    LocalMux I__8686 (
            .O(N__35285),
            .I(\processor_zipi8.arith_logical_result_4 ));
    Odrv4 I__8685 (
            .O(N__35280),
            .I(\processor_zipi8.arith_logical_result_4 ));
    Odrv12 I__8684 (
            .O(N__35275),
            .I(\processor_zipi8.arith_logical_result_4 ));
    Odrv4 I__8683 (
            .O(N__35268),
            .I(\processor_zipi8.arith_logical_result_4 ));
    Odrv4 I__8682 (
            .O(N__35265),
            .I(\processor_zipi8.arith_logical_result_4 ));
    LocalMux I__8681 (
            .O(N__35262),
            .I(\processor_zipi8.arith_logical_result_4 ));
    Odrv12 I__8680 (
            .O(N__35255),
            .I(\processor_zipi8.arith_logical_result_4 ));
    InMux I__8679 (
            .O(N__35240),
            .I(N__35237));
    LocalMux I__8678 (
            .O(N__35237),
            .I(N__35225));
    CascadeMux I__8677 (
            .O(N__35236),
            .I(N__35222));
    InMux I__8676 (
            .O(N__35235),
            .I(N__35215));
    CascadeMux I__8675 (
            .O(N__35234),
            .I(N__35212));
    CascadeMux I__8674 (
            .O(N__35233),
            .I(N__35208));
    CascadeMux I__8673 (
            .O(N__35232),
            .I(N__35205));
    CascadeMux I__8672 (
            .O(N__35231),
            .I(N__35200));
    CascadeMux I__8671 (
            .O(N__35230),
            .I(N__35197));
    CascadeMux I__8670 (
            .O(N__35229),
            .I(N__35194));
    InMux I__8669 (
            .O(N__35228),
            .I(N__35186));
    Span4Mux_v I__8668 (
            .O(N__35225),
            .I(N__35183));
    InMux I__8667 (
            .O(N__35222),
            .I(N__35180));
    InMux I__8666 (
            .O(N__35221),
            .I(N__35177));
    InMux I__8665 (
            .O(N__35220),
            .I(N__35174));
    CascadeMux I__8664 (
            .O(N__35219),
            .I(N__35171));
    CascadeMux I__8663 (
            .O(N__35218),
            .I(N__35166));
    LocalMux I__8662 (
            .O(N__35215),
            .I(N__35163));
    InMux I__8661 (
            .O(N__35212),
            .I(N__35160));
    CascadeMux I__8660 (
            .O(N__35211),
            .I(N__35157));
    InMux I__8659 (
            .O(N__35208),
            .I(N__35152));
    InMux I__8658 (
            .O(N__35205),
            .I(N__35149));
    CascadeMux I__8657 (
            .O(N__35204),
            .I(N__35146));
    InMux I__8656 (
            .O(N__35203),
            .I(N__35142));
    InMux I__8655 (
            .O(N__35200),
            .I(N__35139));
    InMux I__8654 (
            .O(N__35197),
            .I(N__35136));
    InMux I__8653 (
            .O(N__35194),
            .I(N__35133));
    InMux I__8652 (
            .O(N__35193),
            .I(N__35130));
    CascadeMux I__8651 (
            .O(N__35192),
            .I(N__35127));
    CascadeMux I__8650 (
            .O(N__35191),
            .I(N__35124));
    InMux I__8649 (
            .O(N__35190),
            .I(N__35120));
    InMux I__8648 (
            .O(N__35189),
            .I(N__35117));
    LocalMux I__8647 (
            .O(N__35186),
            .I(N__35114));
    IoSpan4Mux I__8646 (
            .O(N__35183),
            .I(N__35107));
    LocalMux I__8645 (
            .O(N__35180),
            .I(N__35107));
    LocalMux I__8644 (
            .O(N__35177),
            .I(N__35107));
    LocalMux I__8643 (
            .O(N__35174),
            .I(N__35104));
    InMux I__8642 (
            .O(N__35171),
            .I(N__35101));
    InMux I__8641 (
            .O(N__35170),
            .I(N__35098));
    CascadeMux I__8640 (
            .O(N__35169),
            .I(N__35094));
    InMux I__8639 (
            .O(N__35166),
            .I(N__35090));
    Span4Mux_v I__8638 (
            .O(N__35163),
            .I(N__35085));
    LocalMux I__8637 (
            .O(N__35160),
            .I(N__35085));
    InMux I__8636 (
            .O(N__35157),
            .I(N__35082));
    InMux I__8635 (
            .O(N__35156),
            .I(N__35079));
    InMux I__8634 (
            .O(N__35155),
            .I(N__35076));
    LocalMux I__8633 (
            .O(N__35152),
            .I(N__35073));
    LocalMux I__8632 (
            .O(N__35149),
            .I(N__35070));
    InMux I__8631 (
            .O(N__35146),
            .I(N__35067));
    InMux I__8630 (
            .O(N__35145),
            .I(N__35064));
    LocalMux I__8629 (
            .O(N__35142),
            .I(N__35057));
    LocalMux I__8628 (
            .O(N__35139),
            .I(N__35057));
    LocalMux I__8627 (
            .O(N__35136),
            .I(N__35057));
    LocalMux I__8626 (
            .O(N__35133),
            .I(N__35054));
    LocalMux I__8625 (
            .O(N__35130),
            .I(N__35051));
    InMux I__8624 (
            .O(N__35127),
            .I(N__35048));
    InMux I__8623 (
            .O(N__35124),
            .I(N__35045));
    InMux I__8622 (
            .O(N__35123),
            .I(N__35042));
    LocalMux I__8621 (
            .O(N__35120),
            .I(N__35039));
    LocalMux I__8620 (
            .O(N__35117),
            .I(N__35032));
    Span4Mux_v I__8619 (
            .O(N__35114),
            .I(N__35032));
    Span4Mux_s2_h I__8618 (
            .O(N__35107),
            .I(N__35032));
    Span4Mux_v I__8617 (
            .O(N__35104),
            .I(N__35029));
    LocalMux I__8616 (
            .O(N__35101),
            .I(N__35024));
    LocalMux I__8615 (
            .O(N__35098),
            .I(N__35024));
    CascadeMux I__8614 (
            .O(N__35097),
            .I(N__35021));
    InMux I__8613 (
            .O(N__35094),
            .I(N__35018));
    InMux I__8612 (
            .O(N__35093),
            .I(N__35015));
    LocalMux I__8611 (
            .O(N__35090),
            .I(N__35008));
    Span4Mux_h I__8610 (
            .O(N__35085),
            .I(N__35008));
    LocalMux I__8609 (
            .O(N__35082),
            .I(N__35008));
    LocalMux I__8608 (
            .O(N__35079),
            .I(N__35001));
    LocalMux I__8607 (
            .O(N__35076),
            .I(N__35001));
    Span4Mux_s1_h I__8606 (
            .O(N__35073),
            .I(N__34996));
    Span4Mux_v I__8605 (
            .O(N__35070),
            .I(N__34996));
    LocalMux I__8604 (
            .O(N__35067),
            .I(N__34989));
    LocalMux I__8603 (
            .O(N__35064),
            .I(N__34989));
    Span4Mux_s3_v I__8602 (
            .O(N__35057),
            .I(N__34989));
    Span4Mux_v I__8601 (
            .O(N__35054),
            .I(N__34986));
    Span4Mux_s2_v I__8600 (
            .O(N__35051),
            .I(N__34979));
    LocalMux I__8599 (
            .O(N__35048),
            .I(N__34979));
    LocalMux I__8598 (
            .O(N__35045),
            .I(N__34979));
    LocalMux I__8597 (
            .O(N__35042),
            .I(N__34968));
    Span4Mux_v I__8596 (
            .O(N__35039),
            .I(N__34968));
    Span4Mux_v I__8595 (
            .O(N__35032),
            .I(N__34968));
    Span4Mux_s2_h I__8594 (
            .O(N__35029),
            .I(N__34968));
    Span4Mux_s2_h I__8593 (
            .O(N__35024),
            .I(N__34968));
    InMux I__8592 (
            .O(N__35021),
            .I(N__34965));
    LocalMux I__8591 (
            .O(N__35018),
            .I(N__34960));
    LocalMux I__8590 (
            .O(N__35015),
            .I(N__34960));
    Span4Mux_h I__8589 (
            .O(N__35008),
            .I(N__34957));
    InMux I__8588 (
            .O(N__35007),
            .I(N__34954));
    InMux I__8587 (
            .O(N__35006),
            .I(N__34951));
    Span12Mux_s8_v I__8586 (
            .O(N__35001),
            .I(N__34948));
    Span4Mux_h I__8585 (
            .O(N__34996),
            .I(N__34945));
    Span4Mux_v I__8584 (
            .O(N__34989),
            .I(N__34940));
    Span4Mux_v I__8583 (
            .O(N__34986),
            .I(N__34940));
    Span4Mux_v I__8582 (
            .O(N__34979),
            .I(N__34935));
    Span4Mux_h I__8581 (
            .O(N__34968),
            .I(N__34935));
    LocalMux I__8580 (
            .O(N__34965),
            .I(N__34926));
    Span12Mux_s6_h I__8579 (
            .O(N__34960),
            .I(N__34926));
    Sp12to4 I__8578 (
            .O(N__34957),
            .I(N__34926));
    LocalMux I__8577 (
            .O(N__34954),
            .I(N__34926));
    LocalMux I__8576 (
            .O(N__34951),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ));
    Odrv12 I__8575 (
            .O(N__34948),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ));
    Odrv4 I__8574 (
            .O(N__34945),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ));
    Odrv4 I__8573 (
            .O(N__34940),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ));
    Odrv4 I__8572 (
            .O(N__34935),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ));
    Odrv12 I__8571 (
            .O(N__34926),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ));
    InMux I__8570 (
            .O(N__34913),
            .I(N__34892));
    InMux I__8569 (
            .O(N__34912),
            .I(N__34892));
    InMux I__8568 (
            .O(N__34911),
            .I(N__34892));
    InMux I__8567 (
            .O(N__34910),
            .I(N__34892));
    InMux I__8566 (
            .O(N__34909),
            .I(N__34892));
    InMux I__8565 (
            .O(N__34908),
            .I(N__34892));
    InMux I__8564 (
            .O(N__34907),
            .I(N__34892));
    LocalMux I__8563 (
            .O(N__34892),
            .I(N__34877));
    InMux I__8562 (
            .O(N__34891),
            .I(N__34862));
    InMux I__8561 (
            .O(N__34890),
            .I(N__34862));
    InMux I__8560 (
            .O(N__34889),
            .I(N__34862));
    InMux I__8559 (
            .O(N__34888),
            .I(N__34862));
    InMux I__8558 (
            .O(N__34887),
            .I(N__34862));
    InMux I__8557 (
            .O(N__34886),
            .I(N__34862));
    InMux I__8556 (
            .O(N__34885),
            .I(N__34862));
    InMux I__8555 (
            .O(N__34884),
            .I(N__34859));
    InMux I__8554 (
            .O(N__34883),
            .I(N__34852));
    InMux I__8553 (
            .O(N__34882),
            .I(N__34852));
    InMux I__8552 (
            .O(N__34881),
            .I(N__34852));
    CascadeMux I__8551 (
            .O(N__34880),
            .I(N__34847));
    Span4Mux_v I__8550 (
            .O(N__34877),
            .I(N__34786));
    LocalMux I__8549 (
            .O(N__34862),
            .I(N__34786));
    LocalMux I__8548 (
            .O(N__34859),
            .I(N__34786));
    LocalMux I__8547 (
            .O(N__34852),
            .I(N__34783));
    InMux I__8546 (
            .O(N__34851),
            .I(N__34766));
    InMux I__8545 (
            .O(N__34850),
            .I(N__34766));
    InMux I__8544 (
            .O(N__34847),
            .I(N__34766));
    InMux I__8543 (
            .O(N__34846),
            .I(N__34766));
    InMux I__8542 (
            .O(N__34845),
            .I(N__34766));
    InMux I__8541 (
            .O(N__34844),
            .I(N__34766));
    InMux I__8540 (
            .O(N__34843),
            .I(N__34766));
    InMux I__8539 (
            .O(N__34842),
            .I(N__34766));
    CascadeMux I__8538 (
            .O(N__34841),
            .I(N__34761));
    CascadeMux I__8537 (
            .O(N__34840),
            .I(N__34757));
    CascadeMux I__8536 (
            .O(N__34839),
            .I(N__34748));
    InMux I__8535 (
            .O(N__34838),
            .I(N__34727));
    InMux I__8534 (
            .O(N__34837),
            .I(N__34727));
    InMux I__8533 (
            .O(N__34836),
            .I(N__34727));
    InMux I__8532 (
            .O(N__34835),
            .I(N__34727));
    InMux I__8531 (
            .O(N__34834),
            .I(N__34727));
    InMux I__8530 (
            .O(N__34833),
            .I(N__34727));
    InMux I__8529 (
            .O(N__34832),
            .I(N__34727));
    InMux I__8528 (
            .O(N__34831),
            .I(N__34723));
    InMux I__8527 (
            .O(N__34830),
            .I(N__34712));
    InMux I__8526 (
            .O(N__34829),
            .I(N__34712));
    InMux I__8525 (
            .O(N__34828),
            .I(N__34712));
    InMux I__8524 (
            .O(N__34827),
            .I(N__34712));
    InMux I__8523 (
            .O(N__34826),
            .I(N__34712));
    CascadeMux I__8522 (
            .O(N__34825),
            .I(N__34708));
    CascadeMux I__8521 (
            .O(N__34824),
            .I(N__34705));
    InMux I__8520 (
            .O(N__34823),
            .I(N__34686));
    InMux I__8519 (
            .O(N__34822),
            .I(N__34686));
    InMux I__8518 (
            .O(N__34821),
            .I(N__34686));
    InMux I__8517 (
            .O(N__34820),
            .I(N__34686));
    InMux I__8516 (
            .O(N__34819),
            .I(N__34686));
    InMux I__8515 (
            .O(N__34818),
            .I(N__34686));
    InMux I__8514 (
            .O(N__34817),
            .I(N__34669));
    InMux I__8513 (
            .O(N__34816),
            .I(N__34669));
    InMux I__8512 (
            .O(N__34815),
            .I(N__34669));
    InMux I__8511 (
            .O(N__34814),
            .I(N__34669));
    InMux I__8510 (
            .O(N__34813),
            .I(N__34669));
    InMux I__8509 (
            .O(N__34812),
            .I(N__34669));
    InMux I__8508 (
            .O(N__34811),
            .I(N__34669));
    InMux I__8507 (
            .O(N__34810),
            .I(N__34669));
    InMux I__8506 (
            .O(N__34809),
            .I(N__34658));
    InMux I__8505 (
            .O(N__34808),
            .I(N__34658));
    InMux I__8504 (
            .O(N__34807),
            .I(N__34658));
    InMux I__8503 (
            .O(N__34806),
            .I(N__34658));
    InMux I__8502 (
            .O(N__34805),
            .I(N__34658));
    InMux I__8501 (
            .O(N__34804),
            .I(N__34640));
    InMux I__8500 (
            .O(N__34803),
            .I(N__34640));
    InMux I__8499 (
            .O(N__34802),
            .I(N__34640));
    InMux I__8498 (
            .O(N__34801),
            .I(N__34640));
    InMux I__8497 (
            .O(N__34800),
            .I(N__34640));
    InMux I__8496 (
            .O(N__34799),
            .I(N__34640));
    InMux I__8495 (
            .O(N__34798),
            .I(N__34626));
    InMux I__8494 (
            .O(N__34797),
            .I(N__34626));
    InMux I__8493 (
            .O(N__34796),
            .I(N__34626));
    CascadeMux I__8492 (
            .O(N__34795),
            .I(N__34621));
    CascadeMux I__8491 (
            .O(N__34794),
            .I(N__34606));
    CascadeMux I__8490 (
            .O(N__34793),
            .I(N__34603));
    Span4Mux_s2_h I__8489 (
            .O(N__34786),
            .I(N__34572));
    Span4Mux_s2_v I__8488 (
            .O(N__34783),
            .I(N__34572));
    LocalMux I__8487 (
            .O(N__34766),
            .I(N__34572));
    InMux I__8486 (
            .O(N__34765),
            .I(N__34564));
    CascadeMux I__8485 (
            .O(N__34764),
            .I(N__34561));
    InMux I__8484 (
            .O(N__34761),
            .I(N__34553));
    InMux I__8483 (
            .O(N__34760),
            .I(N__34536));
    InMux I__8482 (
            .O(N__34757),
            .I(N__34536));
    InMux I__8481 (
            .O(N__34756),
            .I(N__34536));
    InMux I__8480 (
            .O(N__34755),
            .I(N__34536));
    InMux I__8479 (
            .O(N__34754),
            .I(N__34536));
    InMux I__8478 (
            .O(N__34753),
            .I(N__34536));
    InMux I__8477 (
            .O(N__34752),
            .I(N__34536));
    InMux I__8476 (
            .O(N__34751),
            .I(N__34536));
    InMux I__8475 (
            .O(N__34748),
            .I(N__34521));
    InMux I__8474 (
            .O(N__34747),
            .I(N__34521));
    InMux I__8473 (
            .O(N__34746),
            .I(N__34521));
    InMux I__8472 (
            .O(N__34745),
            .I(N__34521));
    InMux I__8471 (
            .O(N__34744),
            .I(N__34521));
    InMux I__8470 (
            .O(N__34743),
            .I(N__34521));
    InMux I__8469 (
            .O(N__34742),
            .I(N__34521));
    LocalMux I__8468 (
            .O(N__34727),
            .I(N__34496));
    InMux I__8467 (
            .O(N__34726),
            .I(N__34491));
    LocalMux I__8466 (
            .O(N__34723),
            .I(N__34488));
    LocalMux I__8465 (
            .O(N__34712),
            .I(N__34485));
    InMux I__8464 (
            .O(N__34711),
            .I(N__34478));
    InMux I__8463 (
            .O(N__34708),
            .I(N__34478));
    InMux I__8462 (
            .O(N__34705),
            .I(N__34478));
    InMux I__8461 (
            .O(N__34704),
            .I(N__34469));
    InMux I__8460 (
            .O(N__34703),
            .I(N__34469));
    InMux I__8459 (
            .O(N__34702),
            .I(N__34469));
    InMux I__8458 (
            .O(N__34701),
            .I(N__34469));
    CascadeMux I__8457 (
            .O(N__34700),
            .I(N__34464));
    InMux I__8456 (
            .O(N__34699),
            .I(N__34461));
    LocalMux I__8455 (
            .O(N__34686),
            .I(N__34454));
    LocalMux I__8454 (
            .O(N__34669),
            .I(N__34454));
    LocalMux I__8453 (
            .O(N__34658),
            .I(N__34454));
    InMux I__8452 (
            .O(N__34657),
            .I(N__34443));
    InMux I__8451 (
            .O(N__34656),
            .I(N__34443));
    InMux I__8450 (
            .O(N__34655),
            .I(N__34443));
    InMux I__8449 (
            .O(N__34654),
            .I(N__34443));
    InMux I__8448 (
            .O(N__34653),
            .I(N__34443));
    LocalMux I__8447 (
            .O(N__34640),
            .I(N__34440));
    InMux I__8446 (
            .O(N__34639),
            .I(N__34425));
    InMux I__8445 (
            .O(N__34638),
            .I(N__34425));
    InMux I__8444 (
            .O(N__34637),
            .I(N__34425));
    InMux I__8443 (
            .O(N__34636),
            .I(N__34425));
    InMux I__8442 (
            .O(N__34635),
            .I(N__34425));
    InMux I__8441 (
            .O(N__34634),
            .I(N__34425));
    InMux I__8440 (
            .O(N__34633),
            .I(N__34425));
    LocalMux I__8439 (
            .O(N__34626),
            .I(N__34422));
    InMux I__8438 (
            .O(N__34625),
            .I(N__34409));
    InMux I__8437 (
            .O(N__34624),
            .I(N__34409));
    InMux I__8436 (
            .O(N__34621),
            .I(N__34409));
    InMux I__8435 (
            .O(N__34620),
            .I(N__34409));
    InMux I__8434 (
            .O(N__34619),
            .I(N__34409));
    InMux I__8433 (
            .O(N__34618),
            .I(N__34409));
    InMux I__8432 (
            .O(N__34617),
            .I(N__34385));
    InMux I__8431 (
            .O(N__34616),
            .I(N__34385));
    InMux I__8430 (
            .O(N__34615),
            .I(N__34385));
    InMux I__8429 (
            .O(N__34614),
            .I(N__34385));
    InMux I__8428 (
            .O(N__34613),
            .I(N__34385));
    InMux I__8427 (
            .O(N__34612),
            .I(N__34385));
    InMux I__8426 (
            .O(N__34611),
            .I(N__34385));
    InMux I__8425 (
            .O(N__34610),
            .I(N__34385));
    InMux I__8424 (
            .O(N__34609),
            .I(N__34368));
    InMux I__8423 (
            .O(N__34606),
            .I(N__34368));
    InMux I__8422 (
            .O(N__34603),
            .I(N__34368));
    InMux I__8421 (
            .O(N__34602),
            .I(N__34368));
    InMux I__8420 (
            .O(N__34601),
            .I(N__34368));
    InMux I__8419 (
            .O(N__34600),
            .I(N__34368));
    InMux I__8418 (
            .O(N__34599),
            .I(N__34368));
    InMux I__8417 (
            .O(N__34598),
            .I(N__34368));
    InMux I__8416 (
            .O(N__34597),
            .I(N__34351));
    InMux I__8415 (
            .O(N__34596),
            .I(N__34351));
    InMux I__8414 (
            .O(N__34595),
            .I(N__34351));
    InMux I__8413 (
            .O(N__34594),
            .I(N__34351));
    InMux I__8412 (
            .O(N__34593),
            .I(N__34351));
    InMux I__8411 (
            .O(N__34592),
            .I(N__34351));
    InMux I__8410 (
            .O(N__34591),
            .I(N__34351));
    InMux I__8409 (
            .O(N__34590),
            .I(N__34351));
    InMux I__8408 (
            .O(N__34589),
            .I(N__34334));
    InMux I__8407 (
            .O(N__34588),
            .I(N__34334));
    InMux I__8406 (
            .O(N__34587),
            .I(N__34334));
    InMux I__8405 (
            .O(N__34586),
            .I(N__34334));
    InMux I__8404 (
            .O(N__34585),
            .I(N__34334));
    InMux I__8403 (
            .O(N__34584),
            .I(N__34334));
    InMux I__8402 (
            .O(N__34583),
            .I(N__34334));
    InMux I__8401 (
            .O(N__34582),
            .I(N__34334));
    InMux I__8400 (
            .O(N__34581),
            .I(N__34327));
    InMux I__8399 (
            .O(N__34580),
            .I(N__34327));
    InMux I__8398 (
            .O(N__34579),
            .I(N__34327));
    Span4Mux_v I__8397 (
            .O(N__34572),
            .I(N__34322));
    InMux I__8396 (
            .O(N__34571),
            .I(N__34319));
    InMux I__8395 (
            .O(N__34570),
            .I(N__34316));
    InMux I__8394 (
            .O(N__34569),
            .I(N__34313));
    InMux I__8393 (
            .O(N__34568),
            .I(N__34310));
    InMux I__8392 (
            .O(N__34567),
            .I(N__34307));
    LocalMux I__8391 (
            .O(N__34564),
            .I(N__34300));
    InMux I__8390 (
            .O(N__34561),
            .I(N__34287));
    InMux I__8389 (
            .O(N__34560),
            .I(N__34287));
    InMux I__8388 (
            .O(N__34559),
            .I(N__34287));
    InMux I__8387 (
            .O(N__34558),
            .I(N__34287));
    InMux I__8386 (
            .O(N__34557),
            .I(N__34287));
    InMux I__8385 (
            .O(N__34556),
            .I(N__34287));
    LocalMux I__8384 (
            .O(N__34553),
            .I(N__34280));
    LocalMux I__8383 (
            .O(N__34536),
            .I(N__34280));
    LocalMux I__8382 (
            .O(N__34521),
            .I(N__34280));
    InMux I__8381 (
            .O(N__34520),
            .I(N__34277));
    InMux I__8380 (
            .O(N__34519),
            .I(N__34267));
    InMux I__8379 (
            .O(N__34518),
            .I(N__34267));
    InMux I__8378 (
            .O(N__34517),
            .I(N__34267));
    InMux I__8377 (
            .O(N__34516),
            .I(N__34267));
    InMux I__8376 (
            .O(N__34515),
            .I(N__34264));
    InMux I__8375 (
            .O(N__34514),
            .I(N__34247));
    InMux I__8374 (
            .O(N__34513),
            .I(N__34247));
    InMux I__8373 (
            .O(N__34512),
            .I(N__34247));
    InMux I__8372 (
            .O(N__34511),
            .I(N__34247));
    InMux I__8371 (
            .O(N__34510),
            .I(N__34247));
    InMux I__8370 (
            .O(N__34509),
            .I(N__34247));
    InMux I__8369 (
            .O(N__34508),
            .I(N__34247));
    InMux I__8368 (
            .O(N__34507),
            .I(N__34247));
    InMux I__8367 (
            .O(N__34506),
            .I(N__34230));
    InMux I__8366 (
            .O(N__34505),
            .I(N__34230));
    InMux I__8365 (
            .O(N__34504),
            .I(N__34230));
    InMux I__8364 (
            .O(N__34503),
            .I(N__34230));
    InMux I__8363 (
            .O(N__34502),
            .I(N__34230));
    InMux I__8362 (
            .O(N__34501),
            .I(N__34230));
    InMux I__8361 (
            .O(N__34500),
            .I(N__34230));
    InMux I__8360 (
            .O(N__34499),
            .I(N__34230));
    Span4Mux_s3_h I__8359 (
            .O(N__34496),
            .I(N__34227));
    InMux I__8358 (
            .O(N__34495),
            .I(N__34222));
    InMux I__8357 (
            .O(N__34494),
            .I(N__34222));
    LocalMux I__8356 (
            .O(N__34491),
            .I(N__34219));
    Span4Mux_v I__8355 (
            .O(N__34488),
            .I(N__34216));
    Span4Mux_v I__8354 (
            .O(N__34485),
            .I(N__34211));
    LocalMux I__8353 (
            .O(N__34478),
            .I(N__34211));
    LocalMux I__8352 (
            .O(N__34469),
            .I(N__34208));
    CascadeMux I__8351 (
            .O(N__34468),
            .I(N__34184));
    InMux I__8350 (
            .O(N__34467),
            .I(N__34177));
    InMux I__8349 (
            .O(N__34464),
            .I(N__34174));
    LocalMux I__8348 (
            .O(N__34461),
            .I(N__34167));
    Span4Mux_v I__8347 (
            .O(N__34454),
            .I(N__34167));
    LocalMux I__8346 (
            .O(N__34443),
            .I(N__34167));
    Span4Mux_h I__8345 (
            .O(N__34440),
            .I(N__34158));
    LocalMux I__8344 (
            .O(N__34425),
            .I(N__34158));
    Span4Mux_s3_v I__8343 (
            .O(N__34422),
            .I(N__34158));
    LocalMux I__8342 (
            .O(N__34409),
            .I(N__34158));
    InMux I__8341 (
            .O(N__34408),
            .I(N__34143));
    InMux I__8340 (
            .O(N__34407),
            .I(N__34143));
    InMux I__8339 (
            .O(N__34406),
            .I(N__34143));
    InMux I__8338 (
            .O(N__34405),
            .I(N__34143));
    InMux I__8337 (
            .O(N__34404),
            .I(N__34143));
    InMux I__8336 (
            .O(N__34403),
            .I(N__34143));
    InMux I__8335 (
            .O(N__34402),
            .I(N__34143));
    LocalMux I__8334 (
            .O(N__34385),
            .I(N__34134));
    LocalMux I__8333 (
            .O(N__34368),
            .I(N__34134));
    LocalMux I__8332 (
            .O(N__34351),
            .I(N__34134));
    LocalMux I__8331 (
            .O(N__34334),
            .I(N__34134));
    LocalMux I__8330 (
            .O(N__34327),
            .I(N__34131));
    InMux I__8329 (
            .O(N__34326),
            .I(N__34124));
    InMux I__8328 (
            .O(N__34325),
            .I(N__34121));
    Span4Mux_h I__8327 (
            .O(N__34322),
            .I(N__34108));
    LocalMux I__8326 (
            .O(N__34319),
            .I(N__34108));
    LocalMux I__8325 (
            .O(N__34316),
            .I(N__34108));
    LocalMux I__8324 (
            .O(N__34313),
            .I(N__34108));
    LocalMux I__8323 (
            .O(N__34310),
            .I(N__34108));
    LocalMux I__8322 (
            .O(N__34307),
            .I(N__34108));
    InMux I__8321 (
            .O(N__34306),
            .I(N__34105));
    InMux I__8320 (
            .O(N__34305),
            .I(N__34102));
    InMux I__8319 (
            .O(N__34304),
            .I(N__34097));
    InMux I__8318 (
            .O(N__34303),
            .I(N__34097));
    Span4Mux_s2_v I__8317 (
            .O(N__34300),
            .I(N__34092));
    LocalMux I__8316 (
            .O(N__34287),
            .I(N__34092));
    Span4Mux_v I__8315 (
            .O(N__34280),
            .I(N__34089));
    LocalMux I__8314 (
            .O(N__34277),
            .I(N__34086));
    CascadeMux I__8313 (
            .O(N__34276),
            .I(N__34075));
    LocalMux I__8312 (
            .O(N__34267),
            .I(N__34059));
    LocalMux I__8311 (
            .O(N__34264),
            .I(N__34059));
    LocalMux I__8310 (
            .O(N__34247),
            .I(N__34059));
    LocalMux I__8309 (
            .O(N__34230),
            .I(N__34059));
    Span4Mux_v I__8308 (
            .O(N__34227),
            .I(N__34054));
    LocalMux I__8307 (
            .O(N__34222),
            .I(N__34054));
    Span4Mux_v I__8306 (
            .O(N__34219),
            .I(N__34045));
    Span4Mux_s0_h I__8305 (
            .O(N__34216),
            .I(N__34045));
    Span4Mux_v I__8304 (
            .O(N__34211),
            .I(N__34045));
    Span4Mux_v I__8303 (
            .O(N__34208),
            .I(N__34045));
    InMux I__8302 (
            .O(N__34207),
            .I(N__34034));
    InMux I__8301 (
            .O(N__34206),
            .I(N__34034));
    InMux I__8300 (
            .O(N__34205),
            .I(N__34034));
    InMux I__8299 (
            .O(N__34204),
            .I(N__34034));
    InMux I__8298 (
            .O(N__34203),
            .I(N__34034));
    InMux I__8297 (
            .O(N__34202),
            .I(N__34023));
    InMux I__8296 (
            .O(N__34201),
            .I(N__34023));
    InMux I__8295 (
            .O(N__34200),
            .I(N__34023));
    InMux I__8294 (
            .O(N__34199),
            .I(N__34023));
    InMux I__8293 (
            .O(N__34198),
            .I(N__34023));
    InMux I__8292 (
            .O(N__34197),
            .I(N__34006));
    InMux I__8291 (
            .O(N__34196),
            .I(N__34006));
    InMux I__8290 (
            .O(N__34195),
            .I(N__34006));
    InMux I__8289 (
            .O(N__34194),
            .I(N__34006));
    InMux I__8288 (
            .O(N__34193),
            .I(N__34006));
    InMux I__8287 (
            .O(N__34192),
            .I(N__34006));
    InMux I__8286 (
            .O(N__34191),
            .I(N__34006));
    InMux I__8285 (
            .O(N__34190),
            .I(N__34006));
    InMux I__8284 (
            .O(N__34189),
            .I(N__34003));
    InMux I__8283 (
            .O(N__34188),
            .I(N__33988));
    InMux I__8282 (
            .O(N__34187),
            .I(N__33988));
    InMux I__8281 (
            .O(N__34184),
            .I(N__33988));
    InMux I__8280 (
            .O(N__34183),
            .I(N__33988));
    InMux I__8279 (
            .O(N__34182),
            .I(N__33988));
    InMux I__8278 (
            .O(N__34181),
            .I(N__33988));
    InMux I__8277 (
            .O(N__34180),
            .I(N__33988));
    LocalMux I__8276 (
            .O(N__34177),
            .I(N__33979));
    LocalMux I__8275 (
            .O(N__34174),
            .I(N__33979));
    Span4Mux_v I__8274 (
            .O(N__34167),
            .I(N__33979));
    Span4Mux_v I__8273 (
            .O(N__34158),
            .I(N__33979));
    LocalMux I__8272 (
            .O(N__34143),
            .I(N__33976));
    Span4Mux_v I__8271 (
            .O(N__34134),
            .I(N__33971));
    Span4Mux_s2_v I__8270 (
            .O(N__34131),
            .I(N__33971));
    InMux I__8269 (
            .O(N__34130),
            .I(N__33968));
    InMux I__8268 (
            .O(N__34129),
            .I(N__33963));
    InMux I__8267 (
            .O(N__34128),
            .I(N__33963));
    InMux I__8266 (
            .O(N__34127),
            .I(N__33960));
    LocalMux I__8265 (
            .O(N__34124),
            .I(N__33955));
    LocalMux I__8264 (
            .O(N__34121),
            .I(N__33955));
    Span4Mux_s2_v I__8263 (
            .O(N__34108),
            .I(N__33932));
    LocalMux I__8262 (
            .O(N__34105),
            .I(N__33932));
    LocalMux I__8261 (
            .O(N__34102),
            .I(N__33932));
    LocalMux I__8260 (
            .O(N__34097),
            .I(N__33932));
    Span4Mux_v I__8259 (
            .O(N__34092),
            .I(N__33932));
    Span4Mux_s1_h I__8258 (
            .O(N__34089),
            .I(N__33932));
    Span4Mux_s2_v I__8257 (
            .O(N__34086),
            .I(N__33932));
    InMux I__8256 (
            .O(N__34085),
            .I(N__33921));
    InMux I__8255 (
            .O(N__34084),
            .I(N__33921));
    InMux I__8254 (
            .O(N__34083),
            .I(N__33914));
    InMux I__8253 (
            .O(N__34082),
            .I(N__33914));
    InMux I__8252 (
            .O(N__34081),
            .I(N__33914));
    InMux I__8251 (
            .O(N__34080),
            .I(N__33909));
    InMux I__8250 (
            .O(N__34079),
            .I(N__33909));
    CascadeMux I__8249 (
            .O(N__34078),
            .I(N__33905));
    InMux I__8248 (
            .O(N__34075),
            .I(N__33899));
    InMux I__8247 (
            .O(N__34074),
            .I(N__33884));
    InMux I__8246 (
            .O(N__34073),
            .I(N__33884));
    InMux I__8245 (
            .O(N__34072),
            .I(N__33884));
    InMux I__8244 (
            .O(N__34071),
            .I(N__33884));
    InMux I__8243 (
            .O(N__34070),
            .I(N__33884));
    InMux I__8242 (
            .O(N__34069),
            .I(N__33884));
    InMux I__8241 (
            .O(N__34068),
            .I(N__33884));
    Span4Mux_v I__8240 (
            .O(N__34059),
            .I(N__33879));
    Span4Mux_h I__8239 (
            .O(N__34054),
            .I(N__33879));
    Sp12to4 I__8238 (
            .O(N__34045),
            .I(N__33870));
    LocalMux I__8237 (
            .O(N__34034),
            .I(N__33870));
    LocalMux I__8236 (
            .O(N__34023),
            .I(N__33870));
    LocalMux I__8235 (
            .O(N__34006),
            .I(N__33870));
    LocalMux I__8234 (
            .O(N__34003),
            .I(N__33866));
    LocalMux I__8233 (
            .O(N__33988),
            .I(N__33863));
    Span4Mux_h I__8232 (
            .O(N__33979),
            .I(N__33858));
    Span4Mux_h I__8231 (
            .O(N__33976),
            .I(N__33858));
    Sp12to4 I__8230 (
            .O(N__33971),
            .I(N__33855));
    LocalMux I__8229 (
            .O(N__33968),
            .I(N__33846));
    LocalMux I__8228 (
            .O(N__33963),
            .I(N__33846));
    LocalMux I__8227 (
            .O(N__33960),
            .I(N__33846));
    Span4Mux_h I__8226 (
            .O(N__33955),
            .I(N__33846));
    InMux I__8225 (
            .O(N__33954),
            .I(N__33829));
    InMux I__8224 (
            .O(N__33953),
            .I(N__33829));
    InMux I__8223 (
            .O(N__33952),
            .I(N__33829));
    InMux I__8222 (
            .O(N__33951),
            .I(N__33829));
    InMux I__8221 (
            .O(N__33950),
            .I(N__33829));
    InMux I__8220 (
            .O(N__33949),
            .I(N__33829));
    InMux I__8219 (
            .O(N__33948),
            .I(N__33829));
    InMux I__8218 (
            .O(N__33947),
            .I(N__33829));
    Sp12to4 I__8217 (
            .O(N__33932),
            .I(N__33826));
    InMux I__8216 (
            .O(N__33931),
            .I(N__33810));
    InMux I__8215 (
            .O(N__33930),
            .I(N__33810));
    InMux I__8214 (
            .O(N__33929),
            .I(N__33810));
    InMux I__8213 (
            .O(N__33928),
            .I(N__33810));
    InMux I__8212 (
            .O(N__33927),
            .I(N__33810));
    InMux I__8211 (
            .O(N__33926),
            .I(N__33810));
    LocalMux I__8210 (
            .O(N__33921),
            .I(N__33803));
    LocalMux I__8209 (
            .O(N__33914),
            .I(N__33803));
    LocalMux I__8208 (
            .O(N__33909),
            .I(N__33803));
    InMux I__8207 (
            .O(N__33908),
            .I(N__33792));
    InMux I__8206 (
            .O(N__33905),
            .I(N__33792));
    InMux I__8205 (
            .O(N__33904),
            .I(N__33792));
    InMux I__8204 (
            .O(N__33903),
            .I(N__33792));
    InMux I__8203 (
            .O(N__33902),
            .I(N__33792));
    LocalMux I__8202 (
            .O(N__33899),
            .I(N__33787));
    LocalMux I__8201 (
            .O(N__33884),
            .I(N__33787));
    Sp12to4 I__8200 (
            .O(N__33879),
            .I(N__33782));
    Span12Mux_s7_h I__8199 (
            .O(N__33870),
            .I(N__33782));
    InMux I__8198 (
            .O(N__33869),
            .I(N__33779));
    Span4Mux_h I__8197 (
            .O(N__33866),
            .I(N__33772));
    Span4Mux_h I__8196 (
            .O(N__33863),
            .I(N__33772));
    Span4Mux_v I__8195 (
            .O(N__33858),
            .I(N__33772));
    Span12Mux_s7_h I__8194 (
            .O(N__33855),
            .I(N__33763));
    Sp12to4 I__8193 (
            .O(N__33846),
            .I(N__33763));
    LocalMux I__8192 (
            .O(N__33829),
            .I(N__33763));
    Span12Mux_s4_h I__8191 (
            .O(N__33826),
            .I(N__33763));
    InMux I__8190 (
            .O(N__33825),
            .I(N__33760));
    InMux I__8189 (
            .O(N__33824),
            .I(N__33755));
    InMux I__8188 (
            .O(N__33823),
            .I(N__33755));
    LocalMux I__8187 (
            .O(N__33810),
            .I(N__33750));
    Span12Mux_v I__8186 (
            .O(N__33803),
            .I(N__33750));
    LocalMux I__8185 (
            .O(N__33792),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    Odrv4 I__8184 (
            .O(N__33787),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    Odrv12 I__8183 (
            .O(N__33782),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    LocalMux I__8182 (
            .O(N__33779),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    Odrv4 I__8181 (
            .O(N__33772),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    Odrv12 I__8180 (
            .O(N__33763),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    LocalMux I__8179 (
            .O(N__33760),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    LocalMux I__8178 (
            .O(N__33755),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    Odrv12 I__8177 (
            .O(N__33750),
            .I(\processor_zipi8.alu_mux_sel_0 ));
    InMux I__8176 (
            .O(N__33731),
            .I(N__33727));
    InMux I__8175 (
            .O(N__33730),
            .I(N__33724));
    LocalMux I__8174 (
            .O(N__33727),
            .I(N__33719));
    LocalMux I__8173 (
            .O(N__33724),
            .I(N__33719));
    Span4Mux_h I__8172 (
            .O(N__33719),
            .I(N__33716));
    Span4Mux_h I__8171 (
            .O(N__33716),
            .I(N__33713));
    Odrv4 I__8170 (
            .O(N__33713),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_4 ));
    ClkMux I__8169 (
            .O(N__33710),
            .I(N__33395));
    ClkMux I__8168 (
            .O(N__33709),
            .I(N__33395));
    ClkMux I__8167 (
            .O(N__33708),
            .I(N__33395));
    ClkMux I__8166 (
            .O(N__33707),
            .I(N__33395));
    ClkMux I__8165 (
            .O(N__33706),
            .I(N__33395));
    ClkMux I__8164 (
            .O(N__33705),
            .I(N__33395));
    ClkMux I__8163 (
            .O(N__33704),
            .I(N__33395));
    ClkMux I__8162 (
            .O(N__33703),
            .I(N__33395));
    ClkMux I__8161 (
            .O(N__33702),
            .I(N__33395));
    ClkMux I__8160 (
            .O(N__33701),
            .I(N__33395));
    ClkMux I__8159 (
            .O(N__33700),
            .I(N__33395));
    ClkMux I__8158 (
            .O(N__33699),
            .I(N__33395));
    ClkMux I__8157 (
            .O(N__33698),
            .I(N__33395));
    ClkMux I__8156 (
            .O(N__33697),
            .I(N__33395));
    ClkMux I__8155 (
            .O(N__33696),
            .I(N__33395));
    ClkMux I__8154 (
            .O(N__33695),
            .I(N__33395));
    ClkMux I__8153 (
            .O(N__33694),
            .I(N__33395));
    ClkMux I__8152 (
            .O(N__33693),
            .I(N__33395));
    ClkMux I__8151 (
            .O(N__33692),
            .I(N__33395));
    ClkMux I__8150 (
            .O(N__33691),
            .I(N__33395));
    ClkMux I__8149 (
            .O(N__33690),
            .I(N__33395));
    ClkMux I__8148 (
            .O(N__33689),
            .I(N__33395));
    ClkMux I__8147 (
            .O(N__33688),
            .I(N__33395));
    ClkMux I__8146 (
            .O(N__33687),
            .I(N__33395));
    ClkMux I__8145 (
            .O(N__33686),
            .I(N__33395));
    ClkMux I__8144 (
            .O(N__33685),
            .I(N__33395));
    ClkMux I__8143 (
            .O(N__33684),
            .I(N__33395));
    ClkMux I__8142 (
            .O(N__33683),
            .I(N__33395));
    ClkMux I__8141 (
            .O(N__33682),
            .I(N__33395));
    ClkMux I__8140 (
            .O(N__33681),
            .I(N__33395));
    ClkMux I__8139 (
            .O(N__33680),
            .I(N__33395));
    ClkMux I__8138 (
            .O(N__33679),
            .I(N__33395));
    ClkMux I__8137 (
            .O(N__33678),
            .I(N__33395));
    ClkMux I__8136 (
            .O(N__33677),
            .I(N__33395));
    ClkMux I__8135 (
            .O(N__33676),
            .I(N__33395));
    ClkMux I__8134 (
            .O(N__33675),
            .I(N__33395));
    ClkMux I__8133 (
            .O(N__33674),
            .I(N__33395));
    ClkMux I__8132 (
            .O(N__33673),
            .I(N__33395));
    ClkMux I__8131 (
            .O(N__33672),
            .I(N__33395));
    ClkMux I__8130 (
            .O(N__33671),
            .I(N__33395));
    ClkMux I__8129 (
            .O(N__33670),
            .I(N__33395));
    ClkMux I__8128 (
            .O(N__33669),
            .I(N__33395));
    ClkMux I__8127 (
            .O(N__33668),
            .I(N__33395));
    ClkMux I__8126 (
            .O(N__33667),
            .I(N__33395));
    ClkMux I__8125 (
            .O(N__33666),
            .I(N__33395));
    ClkMux I__8124 (
            .O(N__33665),
            .I(N__33395));
    ClkMux I__8123 (
            .O(N__33664),
            .I(N__33395));
    ClkMux I__8122 (
            .O(N__33663),
            .I(N__33395));
    ClkMux I__8121 (
            .O(N__33662),
            .I(N__33395));
    ClkMux I__8120 (
            .O(N__33661),
            .I(N__33395));
    ClkMux I__8119 (
            .O(N__33660),
            .I(N__33395));
    ClkMux I__8118 (
            .O(N__33659),
            .I(N__33395));
    ClkMux I__8117 (
            .O(N__33658),
            .I(N__33395));
    ClkMux I__8116 (
            .O(N__33657),
            .I(N__33395));
    ClkMux I__8115 (
            .O(N__33656),
            .I(N__33395));
    ClkMux I__8114 (
            .O(N__33655),
            .I(N__33395));
    ClkMux I__8113 (
            .O(N__33654),
            .I(N__33395));
    ClkMux I__8112 (
            .O(N__33653),
            .I(N__33395));
    ClkMux I__8111 (
            .O(N__33652),
            .I(N__33395));
    ClkMux I__8110 (
            .O(N__33651),
            .I(N__33395));
    ClkMux I__8109 (
            .O(N__33650),
            .I(N__33395));
    ClkMux I__8108 (
            .O(N__33649),
            .I(N__33395));
    ClkMux I__8107 (
            .O(N__33648),
            .I(N__33395));
    ClkMux I__8106 (
            .O(N__33647),
            .I(N__33395));
    ClkMux I__8105 (
            .O(N__33646),
            .I(N__33395));
    ClkMux I__8104 (
            .O(N__33645),
            .I(N__33395));
    ClkMux I__8103 (
            .O(N__33644),
            .I(N__33395));
    ClkMux I__8102 (
            .O(N__33643),
            .I(N__33395));
    ClkMux I__8101 (
            .O(N__33642),
            .I(N__33395));
    ClkMux I__8100 (
            .O(N__33641),
            .I(N__33395));
    ClkMux I__8099 (
            .O(N__33640),
            .I(N__33395));
    ClkMux I__8098 (
            .O(N__33639),
            .I(N__33395));
    ClkMux I__8097 (
            .O(N__33638),
            .I(N__33395));
    ClkMux I__8096 (
            .O(N__33637),
            .I(N__33395));
    ClkMux I__8095 (
            .O(N__33636),
            .I(N__33395));
    ClkMux I__8094 (
            .O(N__33635),
            .I(N__33395));
    ClkMux I__8093 (
            .O(N__33634),
            .I(N__33395));
    ClkMux I__8092 (
            .O(N__33633),
            .I(N__33395));
    ClkMux I__8091 (
            .O(N__33632),
            .I(N__33395));
    ClkMux I__8090 (
            .O(N__33631),
            .I(N__33395));
    ClkMux I__8089 (
            .O(N__33630),
            .I(N__33395));
    ClkMux I__8088 (
            .O(N__33629),
            .I(N__33395));
    ClkMux I__8087 (
            .O(N__33628),
            .I(N__33395));
    ClkMux I__8086 (
            .O(N__33627),
            .I(N__33395));
    ClkMux I__8085 (
            .O(N__33626),
            .I(N__33395));
    ClkMux I__8084 (
            .O(N__33625),
            .I(N__33395));
    ClkMux I__8083 (
            .O(N__33624),
            .I(N__33395));
    ClkMux I__8082 (
            .O(N__33623),
            .I(N__33395));
    ClkMux I__8081 (
            .O(N__33622),
            .I(N__33395));
    ClkMux I__8080 (
            .O(N__33621),
            .I(N__33395));
    ClkMux I__8079 (
            .O(N__33620),
            .I(N__33395));
    ClkMux I__8078 (
            .O(N__33619),
            .I(N__33395));
    ClkMux I__8077 (
            .O(N__33618),
            .I(N__33395));
    ClkMux I__8076 (
            .O(N__33617),
            .I(N__33395));
    ClkMux I__8075 (
            .O(N__33616),
            .I(N__33395));
    ClkMux I__8074 (
            .O(N__33615),
            .I(N__33395));
    ClkMux I__8073 (
            .O(N__33614),
            .I(N__33395));
    ClkMux I__8072 (
            .O(N__33613),
            .I(N__33395));
    ClkMux I__8071 (
            .O(N__33612),
            .I(N__33395));
    ClkMux I__8070 (
            .O(N__33611),
            .I(N__33395));
    ClkMux I__8069 (
            .O(N__33610),
            .I(N__33395));
    ClkMux I__8068 (
            .O(N__33609),
            .I(N__33395));
    ClkMux I__8067 (
            .O(N__33608),
            .I(N__33395));
    ClkMux I__8066 (
            .O(N__33607),
            .I(N__33395));
    ClkMux I__8065 (
            .O(N__33606),
            .I(N__33395));
    GlobalMux I__8064 (
            .O(N__33395),
            .I(N__33392));
    gio2CtrlBuf I__8063 (
            .O(N__33392),
            .I(CLK_3P3_MHZ_c_g));
    CEMux I__8062 (
            .O(N__33389),
            .I(N__33386));
    LocalMux I__8061 (
            .O(N__33386),
            .I(N__33382));
    CEMux I__8060 (
            .O(N__33385),
            .I(N__33379));
    Span4Mux_s0_h I__8059 (
            .O(N__33382),
            .I(N__33376));
    LocalMux I__8058 (
            .O(N__33379),
            .I(N__33373));
    Span4Mux_h I__8057 (
            .O(N__33376),
            .I(N__33370));
    Span4Mux_s3_v I__8056 (
            .O(N__33373),
            .I(N__33367));
    Span4Mux_v I__8055 (
            .O(N__33370),
            .I(N__33364));
    Odrv4 I__8054 (
            .O(N__33367),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22 ));
    Odrv4 I__8053 (
            .O(N__33364),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22 ));
    CascadeMux I__8052 (
            .O(N__33359),
            .I(N__33355));
    InMux I__8051 (
            .O(N__33358),
            .I(N__33352));
    InMux I__8050 (
            .O(N__33355),
            .I(N__33349));
    LocalMux I__8049 (
            .O(N__33352),
            .I(N__33346));
    LocalMux I__8048 (
            .O(N__33349),
            .I(N__33343));
    Span4Mux_h I__8047 (
            .O(N__33346),
            .I(N__33328));
    Span4Mux_s3_h I__8046 (
            .O(N__33343),
            .I(N__33328));
    CascadeMux I__8045 (
            .O(N__33342),
            .I(N__33324));
    CascadeMux I__8044 (
            .O(N__33341),
            .I(N__33321));
    InMux I__8043 (
            .O(N__33340),
            .I(N__33313));
    InMux I__8042 (
            .O(N__33339),
            .I(N__33306));
    InMux I__8041 (
            .O(N__33338),
            .I(N__33303));
    CascadeMux I__8040 (
            .O(N__33337),
            .I(N__33298));
    CascadeMux I__8039 (
            .O(N__33336),
            .I(N__33295));
    CascadeMux I__8038 (
            .O(N__33335),
            .I(N__33291));
    InMux I__8037 (
            .O(N__33334),
            .I(N__33287));
    InMux I__8036 (
            .O(N__33333),
            .I(N__33284));
    IoSpan4Mux I__8035 (
            .O(N__33328),
            .I(N__33281));
    InMux I__8034 (
            .O(N__33327),
            .I(N__33278));
    InMux I__8033 (
            .O(N__33324),
            .I(N__33275));
    InMux I__8032 (
            .O(N__33321),
            .I(N__33272));
    CascadeMux I__8031 (
            .O(N__33320),
            .I(N__33267));
    InMux I__8030 (
            .O(N__33319),
            .I(N__33263));
    InMux I__8029 (
            .O(N__33318),
            .I(N__33260));
    CascadeMux I__8028 (
            .O(N__33317),
            .I(N__33257));
    InMux I__8027 (
            .O(N__33316),
            .I(N__33253));
    LocalMux I__8026 (
            .O(N__33313),
            .I(N__33250));
    InMux I__8025 (
            .O(N__33312),
            .I(N__33247));
    InMux I__8024 (
            .O(N__33311),
            .I(N__33244));
    InMux I__8023 (
            .O(N__33310),
            .I(N__33241));
    InMux I__8022 (
            .O(N__33309),
            .I(N__33238));
    LocalMux I__8021 (
            .O(N__33306),
            .I(N__33235));
    LocalMux I__8020 (
            .O(N__33303),
            .I(N__33232));
    InMux I__8019 (
            .O(N__33302),
            .I(N__33229));
    InMux I__8018 (
            .O(N__33301),
            .I(N__33226));
    InMux I__8017 (
            .O(N__33298),
            .I(N__33223));
    InMux I__8016 (
            .O(N__33295),
            .I(N__33220));
    CascadeMux I__8015 (
            .O(N__33294),
            .I(N__33216));
    InMux I__8014 (
            .O(N__33291),
            .I(N__33213));
    InMux I__8013 (
            .O(N__33290),
            .I(N__33210));
    LocalMux I__8012 (
            .O(N__33287),
            .I(N__33207));
    LocalMux I__8011 (
            .O(N__33284),
            .I(N__33204));
    Span4Mux_s0_v I__8010 (
            .O(N__33281),
            .I(N__33194));
    LocalMux I__8009 (
            .O(N__33278),
            .I(N__33194));
    LocalMux I__8008 (
            .O(N__33275),
            .I(N__33194));
    LocalMux I__8007 (
            .O(N__33272),
            .I(N__33194));
    InMux I__8006 (
            .O(N__33271),
            .I(N__33191));
    InMux I__8005 (
            .O(N__33270),
            .I(N__33186));
    InMux I__8004 (
            .O(N__33267),
            .I(N__33186));
    InMux I__8003 (
            .O(N__33266),
            .I(N__33183));
    LocalMux I__8002 (
            .O(N__33263),
            .I(N__33178));
    LocalMux I__8001 (
            .O(N__33260),
            .I(N__33178));
    InMux I__8000 (
            .O(N__33257),
            .I(N__33175));
    InMux I__7999 (
            .O(N__33256),
            .I(N__33171));
    LocalMux I__7998 (
            .O(N__33253),
            .I(N__33164));
    Span4Mux_v I__7997 (
            .O(N__33250),
            .I(N__33164));
    LocalMux I__7996 (
            .O(N__33247),
            .I(N__33164));
    LocalMux I__7995 (
            .O(N__33244),
            .I(N__33161));
    LocalMux I__7994 (
            .O(N__33241),
            .I(N__33148));
    LocalMux I__7993 (
            .O(N__33238),
            .I(N__33148));
    Span4Mux_s3_h I__7992 (
            .O(N__33235),
            .I(N__33148));
    Span4Mux_v I__7991 (
            .O(N__33232),
            .I(N__33148));
    LocalMux I__7990 (
            .O(N__33229),
            .I(N__33148));
    LocalMux I__7989 (
            .O(N__33226),
            .I(N__33148));
    LocalMux I__7988 (
            .O(N__33223),
            .I(N__33142));
    LocalMux I__7987 (
            .O(N__33220),
            .I(N__33142));
    InMux I__7986 (
            .O(N__33219),
            .I(N__33139));
    InMux I__7985 (
            .O(N__33216),
            .I(N__33136));
    LocalMux I__7984 (
            .O(N__33213),
            .I(N__33133));
    LocalMux I__7983 (
            .O(N__33210),
            .I(N__33130));
    Span4Mux_v I__7982 (
            .O(N__33207),
            .I(N__33125));
    Span4Mux_s0_h I__7981 (
            .O(N__33204),
            .I(N__33125));
    InMux I__7980 (
            .O(N__33203),
            .I(N__33122));
    Span4Mux_h I__7979 (
            .O(N__33194),
            .I(N__33119));
    LocalMux I__7978 (
            .O(N__33191),
            .I(N__33114));
    LocalMux I__7977 (
            .O(N__33186),
            .I(N__33114));
    LocalMux I__7976 (
            .O(N__33183),
            .I(N__33111));
    Span4Mux_v I__7975 (
            .O(N__33178),
            .I(N__33108));
    LocalMux I__7974 (
            .O(N__33175),
            .I(N__33105));
    InMux I__7973 (
            .O(N__33174),
            .I(N__33102));
    LocalMux I__7972 (
            .O(N__33171),
            .I(N__33093));
    Span4Mux_h I__7971 (
            .O(N__33164),
            .I(N__33093));
    Span4Mux_s1_v I__7970 (
            .O(N__33161),
            .I(N__33093));
    Span4Mux_h I__7969 (
            .O(N__33148),
            .I(N__33093));
    CascadeMux I__7968 (
            .O(N__33147),
            .I(N__33090));
    Span4Mux_v I__7967 (
            .O(N__33142),
            .I(N__33087));
    LocalMux I__7966 (
            .O(N__33139),
            .I(N__33080));
    LocalMux I__7965 (
            .O(N__33136),
            .I(N__33080));
    Span4Mux_s3_v I__7964 (
            .O(N__33133),
            .I(N__33080));
    Span4Mux_v I__7963 (
            .O(N__33130),
            .I(N__33077));
    Span4Mux_h I__7962 (
            .O(N__33125),
            .I(N__33072));
    LocalMux I__7961 (
            .O(N__33122),
            .I(N__33072));
    Span4Mux_v I__7960 (
            .O(N__33119),
            .I(N__33067));
    Span4Mux_s3_h I__7959 (
            .O(N__33114),
            .I(N__33067));
    Span4Mux_v I__7958 (
            .O(N__33111),
            .I(N__33062));
    Span4Mux_s1_h I__7957 (
            .O(N__33108),
            .I(N__33062));
    Span12Mux_s7_h I__7956 (
            .O(N__33105),
            .I(N__33059));
    LocalMux I__7955 (
            .O(N__33102),
            .I(N__33054));
    Span4Mux_v I__7954 (
            .O(N__33093),
            .I(N__33054));
    InMux I__7953 (
            .O(N__33090),
            .I(N__33051));
    Span4Mux_h I__7952 (
            .O(N__33087),
            .I(N__33040));
    Span4Mux_v I__7951 (
            .O(N__33080),
            .I(N__33040));
    Span4Mux_h I__7950 (
            .O(N__33077),
            .I(N__33040));
    Span4Mux_v I__7949 (
            .O(N__33072),
            .I(N__33040));
    Span4Mux_v I__7948 (
            .O(N__33067),
            .I(N__33040));
    Odrv4 I__7947 (
            .O(N__33062),
            .I(\processor_zipi8.arith_logical_result_7 ));
    Odrv12 I__7946 (
            .O(N__33059),
            .I(\processor_zipi8.arith_logical_result_7 ));
    Odrv4 I__7945 (
            .O(N__33054),
            .I(\processor_zipi8.arith_logical_result_7 ));
    LocalMux I__7944 (
            .O(N__33051),
            .I(\processor_zipi8.arith_logical_result_7 ));
    Odrv4 I__7943 (
            .O(N__33040),
            .I(\processor_zipi8.arith_logical_result_7 ));
    CascadeMux I__7942 (
            .O(N__33029),
            .I(N__33025));
    CascadeMux I__7941 (
            .O(N__33028),
            .I(N__33022));
    InMux I__7940 (
            .O(N__33025),
            .I(N__33018));
    InMux I__7939 (
            .O(N__33022),
            .I(N__33006));
    CascadeMux I__7938 (
            .O(N__33021),
            .I(N__33003));
    LocalMux I__7937 (
            .O(N__33018),
            .I(N__32996));
    CascadeMux I__7936 (
            .O(N__33017),
            .I(N__32990));
    InMux I__7935 (
            .O(N__33016),
            .I(N__32987));
    InMux I__7934 (
            .O(N__33015),
            .I(N__32984));
    CascadeMux I__7933 (
            .O(N__33014),
            .I(N__32981));
    CascadeMux I__7932 (
            .O(N__33013),
            .I(N__32975));
    CascadeMux I__7931 (
            .O(N__33012),
            .I(N__32970));
    CascadeMux I__7930 (
            .O(N__33011),
            .I(N__32967));
    CascadeMux I__7929 (
            .O(N__33010),
            .I(N__32964));
    CascadeMux I__7928 (
            .O(N__33009),
            .I(N__32961));
    LocalMux I__7927 (
            .O(N__33006),
            .I(N__32957));
    InMux I__7926 (
            .O(N__33003),
            .I(N__32954));
    InMux I__7925 (
            .O(N__33002),
            .I(N__32951));
    CascadeMux I__7924 (
            .O(N__33001),
            .I(N__32948));
    InMux I__7923 (
            .O(N__33000),
            .I(N__32945));
    CascadeMux I__7922 (
            .O(N__32999),
            .I(N__32941));
    Span4Mux_v I__7921 (
            .O(N__32996),
            .I(N__32938));
    CascadeMux I__7920 (
            .O(N__32995),
            .I(N__32935));
    CascadeMux I__7919 (
            .O(N__32994),
            .I(N__32932));
    InMux I__7918 (
            .O(N__32993),
            .I(N__32929));
    InMux I__7917 (
            .O(N__32990),
            .I(N__32926));
    LocalMux I__7916 (
            .O(N__32987),
            .I(N__32923));
    LocalMux I__7915 (
            .O(N__32984),
            .I(N__32920));
    InMux I__7914 (
            .O(N__32981),
            .I(N__32917));
    InMux I__7913 (
            .O(N__32980),
            .I(N__32914));
    InMux I__7912 (
            .O(N__32979),
            .I(N__32911));
    InMux I__7911 (
            .O(N__32978),
            .I(N__32908));
    InMux I__7910 (
            .O(N__32975),
            .I(N__32905));
    InMux I__7909 (
            .O(N__32974),
            .I(N__32902));
    InMux I__7908 (
            .O(N__32973),
            .I(N__32899));
    InMux I__7907 (
            .O(N__32970),
            .I(N__32895));
    InMux I__7906 (
            .O(N__32967),
            .I(N__32892));
    InMux I__7905 (
            .O(N__32964),
            .I(N__32889));
    InMux I__7904 (
            .O(N__32961),
            .I(N__32886));
    CascadeMux I__7903 (
            .O(N__32960),
            .I(N__32883));
    Span4Mux_h I__7902 (
            .O(N__32957),
            .I(N__32876));
    LocalMux I__7901 (
            .O(N__32954),
            .I(N__32876));
    LocalMux I__7900 (
            .O(N__32951),
            .I(N__32876));
    InMux I__7899 (
            .O(N__32948),
            .I(N__32873));
    LocalMux I__7898 (
            .O(N__32945),
            .I(N__32869));
    InMux I__7897 (
            .O(N__32944),
            .I(N__32866));
    InMux I__7896 (
            .O(N__32941),
            .I(N__32863));
    Span4Mux_v I__7895 (
            .O(N__32938),
            .I(N__32860));
    InMux I__7894 (
            .O(N__32935),
            .I(N__32857));
    InMux I__7893 (
            .O(N__32932),
            .I(N__32854));
    LocalMux I__7892 (
            .O(N__32929),
            .I(N__32849));
    LocalMux I__7891 (
            .O(N__32926),
            .I(N__32849));
    Span4Mux_s0_v I__7890 (
            .O(N__32923),
            .I(N__32838));
    Span4Mux_s0_v I__7889 (
            .O(N__32920),
            .I(N__32838));
    LocalMux I__7888 (
            .O(N__32917),
            .I(N__32838));
    LocalMux I__7887 (
            .O(N__32914),
            .I(N__32838));
    LocalMux I__7886 (
            .O(N__32911),
            .I(N__32838));
    LocalMux I__7885 (
            .O(N__32908),
            .I(N__32835));
    LocalMux I__7884 (
            .O(N__32905),
            .I(N__32828));
    LocalMux I__7883 (
            .O(N__32902),
            .I(N__32828));
    LocalMux I__7882 (
            .O(N__32899),
            .I(N__32828));
    CascadeMux I__7881 (
            .O(N__32898),
            .I(N__32825));
    LocalMux I__7880 (
            .O(N__32895),
            .I(N__32820));
    LocalMux I__7879 (
            .O(N__32892),
            .I(N__32817));
    LocalMux I__7878 (
            .O(N__32889),
            .I(N__32812));
    LocalMux I__7877 (
            .O(N__32886),
            .I(N__32812));
    InMux I__7876 (
            .O(N__32883),
            .I(N__32809));
    Span4Mux_s3_v I__7875 (
            .O(N__32876),
            .I(N__32804));
    LocalMux I__7874 (
            .O(N__32873),
            .I(N__32804));
    InMux I__7873 (
            .O(N__32872),
            .I(N__32801));
    Span4Mux_s0_h I__7872 (
            .O(N__32869),
            .I(N__32794));
    LocalMux I__7871 (
            .O(N__32866),
            .I(N__32794));
    LocalMux I__7870 (
            .O(N__32863),
            .I(N__32794));
    Span4Mux_h I__7869 (
            .O(N__32860),
            .I(N__32777));
    LocalMux I__7868 (
            .O(N__32857),
            .I(N__32777));
    LocalMux I__7867 (
            .O(N__32854),
            .I(N__32777));
    Span4Mux_v I__7866 (
            .O(N__32849),
            .I(N__32777));
    Span4Mux_v I__7865 (
            .O(N__32838),
            .I(N__32777));
    Span4Mux_v I__7864 (
            .O(N__32835),
            .I(N__32777));
    Span4Mux_v I__7863 (
            .O(N__32828),
            .I(N__32777));
    InMux I__7862 (
            .O(N__32825),
            .I(N__32772));
    InMux I__7861 (
            .O(N__32824),
            .I(N__32772));
    InMux I__7860 (
            .O(N__32823),
            .I(N__32769));
    Span4Mux_h I__7859 (
            .O(N__32820),
            .I(N__32762));
    Span4Mux_h I__7858 (
            .O(N__32817),
            .I(N__32762));
    Span4Mux_h I__7857 (
            .O(N__32812),
            .I(N__32762));
    LocalMux I__7856 (
            .O(N__32809),
            .I(N__32755));
    Span4Mux_h I__7855 (
            .O(N__32804),
            .I(N__32755));
    LocalMux I__7854 (
            .O(N__32801),
            .I(N__32755));
    Span4Mux_v I__7853 (
            .O(N__32794),
            .I(N__32752));
    InMux I__7852 (
            .O(N__32793),
            .I(N__32749));
    InMux I__7851 (
            .O(N__32792),
            .I(N__32746));
    Sp12to4 I__7850 (
            .O(N__32777),
            .I(N__32741));
    LocalMux I__7849 (
            .O(N__32772),
            .I(N__32741));
    LocalMux I__7848 (
            .O(N__32769),
            .I(N__32736));
    Span4Mux_v I__7847 (
            .O(N__32762),
            .I(N__32736));
    Span4Mux_v I__7846 (
            .O(N__32755),
            .I(N__32733));
    Span4Mux_h I__7845 (
            .O(N__32752),
            .I(N__32730));
    LocalMux I__7844 (
            .O(N__32749),
            .I(N__32723));
    LocalMux I__7843 (
            .O(N__32746),
            .I(N__32723));
    Span12Mux_s7_h I__7842 (
            .O(N__32741),
            .I(N__32723));
    Odrv4 I__7841 (
            .O(N__32736),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269 ));
    Odrv4 I__7840 (
            .O(N__32733),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269 ));
    Odrv4 I__7839 (
            .O(N__32730),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269 ));
    Odrv12 I__7838 (
            .O(N__32723),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269 ));
    CascadeMux I__7837 (
            .O(N__32714),
            .I(N__32711));
    InMux I__7836 (
            .O(N__32711),
            .I(N__32708));
    LocalMux I__7835 (
            .O(N__32708),
            .I(N__32705));
    Span4Mux_s2_v I__7834 (
            .O(N__32705),
            .I(N__32702));
    Span4Mux_v I__7833 (
            .O(N__32702),
            .I(N__32698));
    InMux I__7832 (
            .O(N__32701),
            .I(N__32695));
    Span4Mux_h I__7831 (
            .O(N__32698),
            .I(N__32692));
    LocalMux I__7830 (
            .O(N__32695),
            .I(N__32689));
    Odrv4 I__7829 (
            .O(N__32692),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7 ));
    Odrv12 I__7828 (
            .O(N__32689),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7 ));
    CEMux I__7827 (
            .O(N__32684),
            .I(N__32681));
    LocalMux I__7826 (
            .O(N__32681),
            .I(N__32678));
    Span4Mux_v I__7825 (
            .O(N__32678),
            .I(N__32675));
    IoSpan4Mux I__7824 (
            .O(N__32675),
            .I(N__32671));
    CEMux I__7823 (
            .O(N__32674),
            .I(N__32668));
    IoSpan4Mux I__7822 (
            .O(N__32671),
            .I(N__32665));
    LocalMux I__7821 (
            .O(N__32668),
            .I(N__32662));
    Span4Mux_s2_h I__7820 (
            .O(N__32665),
            .I(N__32659));
    Span12Mux_s3_v I__7819 (
            .O(N__32662),
            .I(N__32656));
    Odrv4 I__7818 (
            .O(N__32659),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21 ));
    Odrv12 I__7817 (
            .O(N__32656),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21 ));
    CascadeMux I__7816 (
            .O(N__32651),
            .I(N__32647));
    CascadeMux I__7815 (
            .O(N__32650),
            .I(N__32644));
    InMux I__7814 (
            .O(N__32647),
            .I(N__32641));
    InMux I__7813 (
            .O(N__32644),
            .I(N__32638));
    LocalMux I__7812 (
            .O(N__32641),
            .I(N__32635));
    LocalMux I__7811 (
            .O(N__32638),
            .I(N__32632));
    Span4Mux_h I__7810 (
            .O(N__32635),
            .I(N__32629));
    Span12Mux_s9_v I__7809 (
            .O(N__32632),
            .I(N__32626));
    Odrv4 I__7808 (
            .O(N__32629),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0 ));
    Odrv12 I__7807 (
            .O(N__32626),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0 ));
    InMux I__7806 (
            .O(N__32621),
            .I(N__32617));
    InMux I__7805 (
            .O(N__32620),
            .I(N__32614));
    LocalMux I__7804 (
            .O(N__32617),
            .I(N__32611));
    LocalMux I__7803 (
            .O(N__32614),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1 ));
    Odrv4 I__7802 (
            .O(N__32611),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1 ));
    InMux I__7801 (
            .O(N__32606),
            .I(N__32602));
    InMux I__7800 (
            .O(N__32605),
            .I(N__32599));
    LocalMux I__7799 (
            .O(N__32602),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1 ));
    LocalMux I__7798 (
            .O(N__32599),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1 ));
    InMux I__7797 (
            .O(N__32594),
            .I(N__32591));
    LocalMux I__7796 (
            .O(N__32591),
            .I(N__32588));
    Odrv12 I__7795 (
            .O(N__32588),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_1 ));
    CascadeMux I__7794 (
            .O(N__32585),
            .I(N__32582));
    InMux I__7793 (
            .O(N__32582),
            .I(N__32578));
    InMux I__7792 (
            .O(N__32581),
            .I(N__32575));
    LocalMux I__7791 (
            .O(N__32578),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2 ));
    LocalMux I__7790 (
            .O(N__32575),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2 ));
    InMux I__7789 (
            .O(N__32570),
            .I(N__32566));
    InMux I__7788 (
            .O(N__32569),
            .I(N__32563));
    LocalMux I__7787 (
            .O(N__32566),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2 ));
    LocalMux I__7786 (
            .O(N__32563),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2 ));
    InMux I__7785 (
            .O(N__32558),
            .I(N__32555));
    LocalMux I__7784 (
            .O(N__32555),
            .I(N__32552));
    Span4Mux_h I__7783 (
            .O(N__32552),
            .I(N__32549));
    Odrv4 I__7782 (
            .O(N__32549),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_2 ));
    CascadeMux I__7781 (
            .O(N__32546),
            .I(N__32542));
    InMux I__7780 (
            .O(N__32545),
            .I(N__32539));
    InMux I__7779 (
            .O(N__32542),
            .I(N__32536));
    LocalMux I__7778 (
            .O(N__32539),
            .I(N__32531));
    LocalMux I__7777 (
            .O(N__32536),
            .I(N__32531));
    Odrv4 I__7776 (
            .O(N__32531),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_3 ));
    CascadeMux I__7775 (
            .O(N__32528),
            .I(N__32525));
    InMux I__7774 (
            .O(N__32525),
            .I(N__32519));
    InMux I__7773 (
            .O(N__32524),
            .I(N__32519));
    LocalMux I__7772 (
            .O(N__32519),
            .I(N__32516));
    Span4Mux_v I__7771 (
            .O(N__32516),
            .I(N__32513));
    Span4Mux_h I__7770 (
            .O(N__32513),
            .I(N__32510));
    Odrv4 I__7769 (
            .O(N__32510),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_4 ));
    CEMux I__7768 (
            .O(N__32507),
            .I(N__32504));
    LocalMux I__7767 (
            .O(N__32504),
            .I(N__32501));
    Span4Mux_s2_h I__7766 (
            .O(N__32501),
            .I(N__32498));
    Span4Mux_h I__7765 (
            .O(N__32498),
            .I(N__32494));
    CEMux I__7764 (
            .O(N__32497),
            .I(N__32491));
    Span4Mux_v I__7763 (
            .O(N__32494),
            .I(N__32488));
    LocalMux I__7762 (
            .O(N__32491),
            .I(N__32485));
    Sp12to4 I__7761 (
            .O(N__32488),
            .I(N__32482));
    Odrv4 I__7760 (
            .O(N__32485),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20 ));
    Odrv12 I__7759 (
            .O(N__32482),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20 ));
    CascadeMux I__7758 (
            .O(N__32477),
            .I(N__32471));
    CascadeMux I__7757 (
            .O(N__32476),
            .I(N__32468));
    CascadeMux I__7756 (
            .O(N__32475),
            .I(N__32465));
    CascadeMux I__7755 (
            .O(N__32474),
            .I(N__32462));
    InMux I__7754 (
            .O(N__32471),
            .I(N__32455));
    InMux I__7753 (
            .O(N__32468),
            .I(N__32452));
    InMux I__7752 (
            .O(N__32465),
            .I(N__32449));
    InMux I__7751 (
            .O(N__32462),
            .I(N__32446));
    InMux I__7750 (
            .O(N__32461),
            .I(N__32443));
    CascadeMux I__7749 (
            .O(N__32460),
            .I(N__32440));
    CascadeMux I__7748 (
            .O(N__32459),
            .I(N__32434));
    CascadeMux I__7747 (
            .O(N__32458),
            .I(N__32428));
    LocalMux I__7746 (
            .O(N__32455),
            .I(N__32423));
    LocalMux I__7745 (
            .O(N__32452),
            .I(N__32423));
    LocalMux I__7744 (
            .O(N__32449),
            .I(N__32416));
    LocalMux I__7743 (
            .O(N__32446),
            .I(N__32416));
    LocalMux I__7742 (
            .O(N__32443),
            .I(N__32416));
    InMux I__7741 (
            .O(N__32440),
            .I(N__32413));
    CascadeMux I__7740 (
            .O(N__32439),
            .I(N__32410));
    InMux I__7739 (
            .O(N__32438),
            .I(N__32407));
    CascadeMux I__7738 (
            .O(N__32437),
            .I(N__32404));
    InMux I__7737 (
            .O(N__32434),
            .I(N__32400));
    CascadeMux I__7736 (
            .O(N__32433),
            .I(N__32395));
    CascadeMux I__7735 (
            .O(N__32432),
            .I(N__32392));
    CascadeMux I__7734 (
            .O(N__32431),
            .I(N__32389));
    InMux I__7733 (
            .O(N__32428),
            .I(N__32386));
    Span4Mux_v I__7732 (
            .O(N__32423),
            .I(N__32381));
    Span4Mux_v I__7731 (
            .O(N__32416),
            .I(N__32381));
    LocalMux I__7730 (
            .O(N__32413),
            .I(N__32377));
    InMux I__7729 (
            .O(N__32410),
            .I(N__32374));
    LocalMux I__7728 (
            .O(N__32407),
            .I(N__32371));
    InMux I__7727 (
            .O(N__32404),
            .I(N__32368));
    CascadeMux I__7726 (
            .O(N__32403),
            .I(N__32365));
    LocalMux I__7725 (
            .O(N__32400),
            .I(N__32359));
    InMux I__7724 (
            .O(N__32399),
            .I(N__32356));
    InMux I__7723 (
            .O(N__32398),
            .I(N__32353));
    InMux I__7722 (
            .O(N__32395),
            .I(N__32346));
    InMux I__7721 (
            .O(N__32392),
            .I(N__32343));
    InMux I__7720 (
            .O(N__32389),
            .I(N__32340));
    LocalMux I__7719 (
            .O(N__32386),
            .I(N__32335));
    IoSpan4Mux I__7718 (
            .O(N__32381),
            .I(N__32335));
    InMux I__7717 (
            .O(N__32380),
            .I(N__32332));
    Span4Mux_h I__7716 (
            .O(N__32377),
            .I(N__32325));
    LocalMux I__7715 (
            .O(N__32374),
            .I(N__32325));
    Span4Mux_s2_h I__7714 (
            .O(N__32371),
            .I(N__32325));
    LocalMux I__7713 (
            .O(N__32368),
            .I(N__32320));
    InMux I__7712 (
            .O(N__32365),
            .I(N__32317));
    CascadeMux I__7711 (
            .O(N__32364),
            .I(N__32313));
    CascadeMux I__7710 (
            .O(N__32363),
            .I(N__32310));
    InMux I__7709 (
            .O(N__32362),
            .I(N__32307));
    Span4Mux_s3_h I__7708 (
            .O(N__32359),
            .I(N__32300));
    LocalMux I__7707 (
            .O(N__32356),
            .I(N__32300));
    LocalMux I__7706 (
            .O(N__32353),
            .I(N__32300));
    CascadeMux I__7705 (
            .O(N__32352),
            .I(N__32296));
    CascadeMux I__7704 (
            .O(N__32351),
            .I(N__32293));
    CascadeMux I__7703 (
            .O(N__32350),
            .I(N__32290));
    InMux I__7702 (
            .O(N__32349),
            .I(N__32286));
    LocalMux I__7701 (
            .O(N__32346),
            .I(N__32279));
    LocalMux I__7700 (
            .O(N__32343),
            .I(N__32279));
    LocalMux I__7699 (
            .O(N__32340),
            .I(N__32279));
    Span4Mux_s2_h I__7698 (
            .O(N__32335),
            .I(N__32276));
    LocalMux I__7697 (
            .O(N__32332),
            .I(N__32271));
    Span4Mux_h I__7696 (
            .O(N__32325),
            .I(N__32271));
    InMux I__7695 (
            .O(N__32324),
            .I(N__32268));
    InMux I__7694 (
            .O(N__32323),
            .I(N__32265));
    Span4Mux_v I__7693 (
            .O(N__32320),
            .I(N__32259));
    LocalMux I__7692 (
            .O(N__32317),
            .I(N__32259));
    CascadeMux I__7691 (
            .O(N__32316),
            .I(N__32256));
    InMux I__7690 (
            .O(N__32313),
            .I(N__32253));
    InMux I__7689 (
            .O(N__32310),
            .I(N__32250));
    LocalMux I__7688 (
            .O(N__32307),
            .I(N__32245));
    Span4Mux_v I__7687 (
            .O(N__32300),
            .I(N__32245));
    CascadeMux I__7686 (
            .O(N__32299),
            .I(N__32241));
    InMux I__7685 (
            .O(N__32296),
            .I(N__32237));
    InMux I__7684 (
            .O(N__32293),
            .I(N__32234));
    InMux I__7683 (
            .O(N__32290),
            .I(N__32231));
    CascadeMux I__7682 (
            .O(N__32289),
            .I(N__32227));
    LocalMux I__7681 (
            .O(N__32286),
            .I(N__32224));
    Span4Mux_v I__7680 (
            .O(N__32279),
            .I(N__32215));
    Span4Mux_h I__7679 (
            .O(N__32276),
            .I(N__32215));
    Span4Mux_v I__7678 (
            .O(N__32271),
            .I(N__32215));
    LocalMux I__7677 (
            .O(N__32268),
            .I(N__32215));
    LocalMux I__7676 (
            .O(N__32265),
            .I(N__32212));
    InMux I__7675 (
            .O(N__32264),
            .I(N__32209));
    Span4Mux_s2_v I__7674 (
            .O(N__32259),
            .I(N__32206));
    InMux I__7673 (
            .O(N__32256),
            .I(N__32203));
    LocalMux I__7672 (
            .O(N__32253),
            .I(N__32200));
    LocalMux I__7671 (
            .O(N__32250),
            .I(N__32195));
    Span4Mux_v I__7670 (
            .O(N__32245),
            .I(N__32195));
    InMux I__7669 (
            .O(N__32244),
            .I(N__32192));
    InMux I__7668 (
            .O(N__32241),
            .I(N__32189));
    InMux I__7667 (
            .O(N__32240),
            .I(N__32186));
    LocalMux I__7666 (
            .O(N__32237),
            .I(N__32179));
    LocalMux I__7665 (
            .O(N__32234),
            .I(N__32179));
    LocalMux I__7664 (
            .O(N__32231),
            .I(N__32179));
    CascadeMux I__7663 (
            .O(N__32230),
            .I(N__32176));
    InMux I__7662 (
            .O(N__32227),
            .I(N__32173));
    Span4Mux_h I__7661 (
            .O(N__32224),
            .I(N__32168));
    Span4Mux_h I__7660 (
            .O(N__32215),
            .I(N__32168));
    Span4Mux_h I__7659 (
            .O(N__32212),
            .I(N__32165));
    LocalMux I__7658 (
            .O(N__32209),
            .I(N__32160));
    Span4Mux_h I__7657 (
            .O(N__32206),
            .I(N__32160));
    LocalMux I__7656 (
            .O(N__32203),
            .I(N__32153));
    Span4Mux_s2_v I__7655 (
            .O(N__32200),
            .I(N__32153));
    Span4Mux_s3_h I__7654 (
            .O(N__32195),
            .I(N__32153));
    LocalMux I__7653 (
            .O(N__32192),
            .I(N__32144));
    LocalMux I__7652 (
            .O(N__32189),
            .I(N__32144));
    LocalMux I__7651 (
            .O(N__32186),
            .I(N__32144));
    Span12Mux_s7_h I__7650 (
            .O(N__32179),
            .I(N__32144));
    InMux I__7649 (
            .O(N__32176),
            .I(N__32141));
    LocalMux I__7648 (
            .O(N__32173),
            .I(N__32136));
    Span4Mux_v I__7647 (
            .O(N__32168),
            .I(N__32136));
    Odrv4 I__7646 (
            .O(N__32165),
            .I(\processor_zipi8.arith_logical_result_0 ));
    Odrv4 I__7645 (
            .O(N__32160),
            .I(\processor_zipi8.arith_logical_result_0 ));
    Odrv4 I__7644 (
            .O(N__32153),
            .I(\processor_zipi8.arith_logical_result_0 ));
    Odrv12 I__7643 (
            .O(N__32144),
            .I(\processor_zipi8.arith_logical_result_0 ));
    LocalMux I__7642 (
            .O(N__32141),
            .I(\processor_zipi8.arith_logical_result_0 ));
    Odrv4 I__7641 (
            .O(N__32136),
            .I(\processor_zipi8.arith_logical_result_0 ));
    InMux I__7640 (
            .O(N__32123),
            .I(N__32116));
    InMux I__7639 (
            .O(N__32122),
            .I(N__32112));
    InMux I__7638 (
            .O(N__32121),
            .I(N__32106));
    InMux I__7637 (
            .O(N__32120),
            .I(N__32103));
    CascadeMux I__7636 (
            .O(N__32119),
            .I(N__32094));
    LocalMux I__7635 (
            .O(N__32116),
            .I(N__32089));
    InMux I__7634 (
            .O(N__32115),
            .I(N__32084));
    LocalMux I__7633 (
            .O(N__32112),
            .I(N__32081));
    CascadeMux I__7632 (
            .O(N__32111),
            .I(N__32076));
    InMux I__7631 (
            .O(N__32110),
            .I(N__32073));
    CascadeMux I__7630 (
            .O(N__32109),
            .I(N__32070));
    LocalMux I__7629 (
            .O(N__32106),
            .I(N__32065));
    LocalMux I__7628 (
            .O(N__32103),
            .I(N__32065));
    InMux I__7627 (
            .O(N__32102),
            .I(N__32062));
    InMux I__7626 (
            .O(N__32101),
            .I(N__32059));
    CascadeMux I__7625 (
            .O(N__32100),
            .I(N__32055));
    CascadeMux I__7624 (
            .O(N__32099),
            .I(N__32052));
    CascadeMux I__7623 (
            .O(N__32098),
            .I(N__32049));
    CascadeMux I__7622 (
            .O(N__32097),
            .I(N__32046));
    InMux I__7621 (
            .O(N__32094),
            .I(N__32043));
    InMux I__7620 (
            .O(N__32093),
            .I(N__32040));
    InMux I__7619 (
            .O(N__32092),
            .I(N__32037));
    Span4Mux_v I__7618 (
            .O(N__32089),
            .I(N__32034));
    InMux I__7617 (
            .O(N__32088),
            .I(N__32031));
    InMux I__7616 (
            .O(N__32087),
            .I(N__32028));
    LocalMux I__7615 (
            .O(N__32084),
            .I(N__32019));
    Span4Mux_s1_h I__7614 (
            .O(N__32081),
            .I(N__32016));
    CascadeMux I__7613 (
            .O(N__32080),
            .I(N__32013));
    InMux I__7612 (
            .O(N__32079),
            .I(N__32010));
    InMux I__7611 (
            .O(N__32076),
            .I(N__32007));
    LocalMux I__7610 (
            .O(N__32073),
            .I(N__32004));
    InMux I__7609 (
            .O(N__32070),
            .I(N__32001));
    Span4Mux_s3_h I__7608 (
            .O(N__32065),
            .I(N__31998));
    LocalMux I__7607 (
            .O(N__32062),
            .I(N__31992));
    LocalMux I__7606 (
            .O(N__32059),
            .I(N__31992));
    InMux I__7605 (
            .O(N__32058),
            .I(N__31989));
    InMux I__7604 (
            .O(N__32055),
            .I(N__31985));
    InMux I__7603 (
            .O(N__32052),
            .I(N__31982));
    InMux I__7602 (
            .O(N__32049),
            .I(N__31979));
    InMux I__7601 (
            .O(N__32046),
            .I(N__31976));
    LocalMux I__7600 (
            .O(N__32043),
            .I(N__31973));
    LocalMux I__7599 (
            .O(N__32040),
            .I(N__31968));
    LocalMux I__7598 (
            .O(N__32037),
            .I(N__31968));
    IoSpan4Mux I__7597 (
            .O(N__32034),
            .I(N__31963));
    LocalMux I__7596 (
            .O(N__32031),
            .I(N__31963));
    LocalMux I__7595 (
            .O(N__32028),
            .I(N__31960));
    CascadeMux I__7594 (
            .O(N__32027),
            .I(N__31955));
    InMux I__7593 (
            .O(N__32026),
            .I(N__31952));
    InMux I__7592 (
            .O(N__32025),
            .I(N__31949));
    InMux I__7591 (
            .O(N__32024),
            .I(N__31946));
    InMux I__7590 (
            .O(N__32023),
            .I(N__31943));
    InMux I__7589 (
            .O(N__32022),
            .I(N__31940));
    Span4Mux_s1_h I__7588 (
            .O(N__32019),
            .I(N__31937));
    Span4Mux_v I__7587 (
            .O(N__32016),
            .I(N__31934));
    InMux I__7586 (
            .O(N__32013),
            .I(N__31931));
    LocalMux I__7585 (
            .O(N__32010),
            .I(N__31920));
    LocalMux I__7584 (
            .O(N__32007),
            .I(N__31920));
    Span4Mux_s3_h I__7583 (
            .O(N__32004),
            .I(N__31920));
    LocalMux I__7582 (
            .O(N__32001),
            .I(N__31920));
    Span4Mux_v I__7581 (
            .O(N__31998),
            .I(N__31920));
    InMux I__7580 (
            .O(N__31997),
            .I(N__31917));
    Span4Mux_s3_h I__7579 (
            .O(N__31992),
            .I(N__31914));
    LocalMux I__7578 (
            .O(N__31989),
            .I(N__31911));
    InMux I__7577 (
            .O(N__31988),
            .I(N__31908));
    LocalMux I__7576 (
            .O(N__31985),
            .I(N__31905));
    LocalMux I__7575 (
            .O(N__31982),
            .I(N__31898));
    LocalMux I__7574 (
            .O(N__31979),
            .I(N__31898));
    LocalMux I__7573 (
            .O(N__31976),
            .I(N__31898));
    Span4Mux_v I__7572 (
            .O(N__31973),
            .I(N__31889));
    Span4Mux_v I__7571 (
            .O(N__31968),
            .I(N__31889));
    Span4Mux_s3_h I__7570 (
            .O(N__31963),
            .I(N__31889));
    Span4Mux_s3_h I__7569 (
            .O(N__31960),
            .I(N__31889));
    InMux I__7568 (
            .O(N__31959),
            .I(N__31886));
    InMux I__7567 (
            .O(N__31958),
            .I(N__31883));
    InMux I__7566 (
            .O(N__31955),
            .I(N__31880));
    LocalMux I__7565 (
            .O(N__31952),
            .I(N__31871));
    LocalMux I__7564 (
            .O(N__31949),
            .I(N__31871));
    LocalMux I__7563 (
            .O(N__31946),
            .I(N__31871));
    LocalMux I__7562 (
            .O(N__31943),
            .I(N__31871));
    LocalMux I__7561 (
            .O(N__31940),
            .I(N__31868));
    Span4Mux_v I__7560 (
            .O(N__31937),
            .I(N__31863));
    Span4Mux_v I__7559 (
            .O(N__31934),
            .I(N__31863));
    LocalMux I__7558 (
            .O(N__31931),
            .I(N__31858));
    Span4Mux_v I__7557 (
            .O(N__31920),
            .I(N__31858));
    LocalMux I__7556 (
            .O(N__31917),
            .I(N__31851));
    Span4Mux_v I__7555 (
            .O(N__31914),
            .I(N__31851));
    Span4Mux_s3_h I__7554 (
            .O(N__31911),
            .I(N__31851));
    LocalMux I__7553 (
            .O(N__31908),
            .I(N__31842));
    Span4Mux_h I__7552 (
            .O(N__31905),
            .I(N__31842));
    Span4Mux_v I__7551 (
            .O(N__31898),
            .I(N__31842));
    Span4Mux_h I__7550 (
            .O(N__31889),
            .I(N__31842));
    LocalMux I__7549 (
            .O(N__31886),
            .I(N__31832));
    LocalMux I__7548 (
            .O(N__31883),
            .I(N__31832));
    LocalMux I__7547 (
            .O(N__31880),
            .I(N__31832));
    Span12Mux_v I__7546 (
            .O(N__31871),
            .I(N__31832));
    Span4Mux_s2_v I__7545 (
            .O(N__31868),
            .I(N__31827));
    Span4Mux_h I__7544 (
            .O(N__31863),
            .I(N__31827));
    Span4Mux_h I__7543 (
            .O(N__31858),
            .I(N__31824));
    Span4Mux_h I__7542 (
            .O(N__31851),
            .I(N__31819));
    Span4Mux_v I__7541 (
            .O(N__31842),
            .I(N__31819));
    InMux I__7540 (
            .O(N__31841),
            .I(N__31816));
    Odrv12 I__7539 (
            .O(N__31832),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197 ));
    Odrv4 I__7538 (
            .O(N__31827),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197 ));
    Odrv4 I__7537 (
            .O(N__31824),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197 ));
    Odrv4 I__7536 (
            .O(N__31819),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197 ));
    LocalMux I__7535 (
            .O(N__31816),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197 ));
    InMux I__7534 (
            .O(N__31805),
            .I(N__31802));
    LocalMux I__7533 (
            .O(N__31802),
            .I(N__31798));
    InMux I__7532 (
            .O(N__31801),
            .I(N__31795));
    Span4Mux_h I__7531 (
            .O(N__31798),
            .I(N__31792));
    LocalMux I__7530 (
            .O(N__31795),
            .I(N__31789));
    Span4Mux_s0_h I__7529 (
            .O(N__31792),
            .I(N__31786));
    Span4Mux_h I__7528 (
            .O(N__31789),
            .I(N__31783));
    Odrv4 I__7527 (
            .O(N__31786),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0 ));
    Odrv4 I__7526 (
            .O(N__31783),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0 ));
    InMux I__7525 (
            .O(N__31778),
            .I(N__31772));
    InMux I__7524 (
            .O(N__31777),
            .I(N__31772));
    LocalMux I__7523 (
            .O(N__31772),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_7 ));
    CascadeMux I__7522 (
            .O(N__31769),
            .I(N__31765));
    InMux I__7521 (
            .O(N__31768),
            .I(N__31760));
    InMux I__7520 (
            .O(N__31765),
            .I(N__31760));
    LocalMux I__7519 (
            .O(N__31760),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_7 ));
    InMux I__7518 (
            .O(N__31757),
            .I(N__31754));
    LocalMux I__7517 (
            .O(N__31754),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_7 ));
    CascadeMux I__7516 (
            .O(N__31751),
            .I(N__31746));
    InMux I__7515 (
            .O(N__31750),
            .I(N__31738));
    InMux I__7514 (
            .O(N__31749),
            .I(N__31725));
    InMux I__7513 (
            .O(N__31746),
            .I(N__31725));
    InMux I__7512 (
            .O(N__31745),
            .I(N__31725));
    InMux I__7511 (
            .O(N__31744),
            .I(N__31722));
    CascadeMux I__7510 (
            .O(N__31743),
            .I(N__31719));
    CascadeMux I__7509 (
            .O(N__31742),
            .I(N__31714));
    CascadeMux I__7508 (
            .O(N__31741),
            .I(N__31709));
    LocalMux I__7507 (
            .O(N__31738),
            .I(N__31685));
    InMux I__7506 (
            .O(N__31737),
            .I(N__31664));
    InMux I__7505 (
            .O(N__31736),
            .I(N__31664));
    InMux I__7504 (
            .O(N__31735),
            .I(N__31664));
    InMux I__7503 (
            .O(N__31734),
            .I(N__31664));
    CascadeMux I__7502 (
            .O(N__31733),
            .I(N__31660));
    CascadeMux I__7501 (
            .O(N__31732),
            .I(N__31657));
    LocalMux I__7500 (
            .O(N__31725),
            .I(N__31652));
    LocalMux I__7499 (
            .O(N__31722),
            .I(N__31652));
    InMux I__7498 (
            .O(N__31719),
            .I(N__31647));
    InMux I__7497 (
            .O(N__31718),
            .I(N__31647));
    InMux I__7496 (
            .O(N__31717),
            .I(N__31642));
    InMux I__7495 (
            .O(N__31714),
            .I(N__31642));
    InMux I__7494 (
            .O(N__31713),
            .I(N__31639));
    InMux I__7493 (
            .O(N__31712),
            .I(N__31632));
    InMux I__7492 (
            .O(N__31709),
            .I(N__31632));
    InMux I__7491 (
            .O(N__31708),
            .I(N__31632));
    InMux I__7490 (
            .O(N__31707),
            .I(N__31625));
    InMux I__7489 (
            .O(N__31706),
            .I(N__31625));
    InMux I__7488 (
            .O(N__31705),
            .I(N__31625));
    CascadeMux I__7487 (
            .O(N__31704),
            .I(N__31620));
    CascadeMux I__7486 (
            .O(N__31703),
            .I(N__31617));
    InMux I__7485 (
            .O(N__31702),
            .I(N__31609));
    InMux I__7484 (
            .O(N__31701),
            .I(N__31606));
    InMux I__7483 (
            .O(N__31700),
            .I(N__31601));
    InMux I__7482 (
            .O(N__31699),
            .I(N__31601));
    InMux I__7481 (
            .O(N__31698),
            .I(N__31598));
    InMux I__7480 (
            .O(N__31697),
            .I(N__31595));
    InMux I__7479 (
            .O(N__31696),
            .I(N__31592));
    CascadeMux I__7478 (
            .O(N__31695),
            .I(N__31586));
    InMux I__7477 (
            .O(N__31694),
            .I(N__31578));
    CascadeMux I__7476 (
            .O(N__31693),
            .I(N__31565));
    InMux I__7475 (
            .O(N__31692),
            .I(N__31558));
    InMux I__7474 (
            .O(N__31691),
            .I(N__31558));
    InMux I__7473 (
            .O(N__31690),
            .I(N__31558));
    InMux I__7472 (
            .O(N__31689),
            .I(N__31553));
    InMux I__7471 (
            .O(N__31688),
            .I(N__31553));
    Span4Mux_h I__7470 (
            .O(N__31685),
            .I(N__31549));
    InMux I__7469 (
            .O(N__31684),
            .I(N__31542));
    InMux I__7468 (
            .O(N__31683),
            .I(N__31542));
    InMux I__7467 (
            .O(N__31682),
            .I(N__31542));
    InMux I__7466 (
            .O(N__31681),
            .I(N__31525));
    InMux I__7465 (
            .O(N__31680),
            .I(N__31525));
    InMux I__7464 (
            .O(N__31679),
            .I(N__31525));
    InMux I__7463 (
            .O(N__31678),
            .I(N__31525));
    InMux I__7462 (
            .O(N__31677),
            .I(N__31525));
    InMux I__7461 (
            .O(N__31676),
            .I(N__31518));
    InMux I__7460 (
            .O(N__31675),
            .I(N__31518));
    InMux I__7459 (
            .O(N__31674),
            .I(N__31518));
    CascadeMux I__7458 (
            .O(N__31673),
            .I(N__31509));
    LocalMux I__7457 (
            .O(N__31664),
            .I(N__31504));
    InMux I__7456 (
            .O(N__31663),
            .I(N__31497));
    InMux I__7455 (
            .O(N__31660),
            .I(N__31497));
    InMux I__7454 (
            .O(N__31657),
            .I(N__31497));
    Span4Mux_v I__7453 (
            .O(N__31652),
            .I(N__31490));
    LocalMux I__7452 (
            .O(N__31647),
            .I(N__31490));
    LocalMux I__7451 (
            .O(N__31642),
            .I(N__31490));
    LocalMux I__7450 (
            .O(N__31639),
            .I(N__31483));
    LocalMux I__7449 (
            .O(N__31632),
            .I(N__31483));
    LocalMux I__7448 (
            .O(N__31625),
            .I(N__31483));
    InMux I__7447 (
            .O(N__31624),
            .I(N__31472));
    InMux I__7446 (
            .O(N__31623),
            .I(N__31472));
    InMux I__7445 (
            .O(N__31620),
            .I(N__31472));
    InMux I__7444 (
            .O(N__31617),
            .I(N__31472));
    InMux I__7443 (
            .O(N__31616),
            .I(N__31472));
    InMux I__7442 (
            .O(N__31615),
            .I(N__31463));
    InMux I__7441 (
            .O(N__31614),
            .I(N__31463));
    InMux I__7440 (
            .O(N__31613),
            .I(N__31463));
    InMux I__7439 (
            .O(N__31612),
            .I(N__31463));
    LocalMux I__7438 (
            .O(N__31609),
            .I(N__31454));
    LocalMux I__7437 (
            .O(N__31606),
            .I(N__31454));
    LocalMux I__7436 (
            .O(N__31601),
            .I(N__31454));
    LocalMux I__7435 (
            .O(N__31598),
            .I(N__31454));
    LocalMux I__7434 (
            .O(N__31595),
            .I(N__31449));
    LocalMux I__7433 (
            .O(N__31592),
            .I(N__31449));
    InMux I__7432 (
            .O(N__31591),
            .I(N__31440));
    InMux I__7431 (
            .O(N__31590),
            .I(N__31440));
    InMux I__7430 (
            .O(N__31589),
            .I(N__31440));
    InMux I__7429 (
            .O(N__31586),
            .I(N__31440));
    InMux I__7428 (
            .O(N__31585),
            .I(N__31429));
    InMux I__7427 (
            .O(N__31584),
            .I(N__31429));
    InMux I__7426 (
            .O(N__31583),
            .I(N__31429));
    InMux I__7425 (
            .O(N__31582),
            .I(N__31429));
    InMux I__7424 (
            .O(N__31581),
            .I(N__31429));
    LocalMux I__7423 (
            .O(N__31578),
            .I(N__31421));
    InMux I__7422 (
            .O(N__31577),
            .I(N__31414));
    InMux I__7421 (
            .O(N__31576),
            .I(N__31414));
    InMux I__7420 (
            .O(N__31575),
            .I(N__31414));
    InMux I__7419 (
            .O(N__31574),
            .I(N__31409));
    InMux I__7418 (
            .O(N__31573),
            .I(N__31409));
    InMux I__7417 (
            .O(N__31572),
            .I(N__31404));
    InMux I__7416 (
            .O(N__31571),
            .I(N__31404));
    InMux I__7415 (
            .O(N__31570),
            .I(N__31399));
    InMux I__7414 (
            .O(N__31569),
            .I(N__31399));
    CascadeMux I__7413 (
            .O(N__31568),
            .I(N__31395));
    InMux I__7412 (
            .O(N__31565),
            .I(N__31387));
    LocalMux I__7411 (
            .O(N__31558),
            .I(N__31381));
    LocalMux I__7410 (
            .O(N__31553),
            .I(N__31378));
    InMux I__7409 (
            .O(N__31552),
            .I(N__31375));
    Span4Mux_h I__7408 (
            .O(N__31549),
            .I(N__31370));
    LocalMux I__7407 (
            .O(N__31542),
            .I(N__31370));
    InMux I__7406 (
            .O(N__31541),
            .I(N__31359));
    InMux I__7405 (
            .O(N__31540),
            .I(N__31359));
    InMux I__7404 (
            .O(N__31539),
            .I(N__31359));
    InMux I__7403 (
            .O(N__31538),
            .I(N__31359));
    InMux I__7402 (
            .O(N__31537),
            .I(N__31359));
    CascadeMux I__7401 (
            .O(N__31536),
            .I(N__31356));
    LocalMux I__7400 (
            .O(N__31525),
            .I(N__31353));
    LocalMux I__7399 (
            .O(N__31518),
            .I(N__31350));
    InMux I__7398 (
            .O(N__31517),
            .I(N__31343));
    InMux I__7397 (
            .O(N__31516),
            .I(N__31343));
    InMux I__7396 (
            .O(N__31515),
            .I(N__31343));
    InMux I__7395 (
            .O(N__31514),
            .I(N__31327));
    InMux I__7394 (
            .O(N__31513),
            .I(N__31327));
    InMux I__7393 (
            .O(N__31512),
            .I(N__31327));
    InMux I__7392 (
            .O(N__31509),
            .I(N__31327));
    CascadeMux I__7391 (
            .O(N__31508),
            .I(N__31322));
    InMux I__7390 (
            .O(N__31507),
            .I(N__31317));
    Span4Mux_v I__7389 (
            .O(N__31504),
            .I(N__31306));
    LocalMux I__7388 (
            .O(N__31497),
            .I(N__31306));
    Span4Mux_h I__7387 (
            .O(N__31490),
            .I(N__31306));
    Span4Mux_v I__7386 (
            .O(N__31483),
            .I(N__31306));
    LocalMux I__7385 (
            .O(N__31472),
            .I(N__31306));
    LocalMux I__7384 (
            .O(N__31463),
            .I(N__31302));
    Span4Mux_v I__7383 (
            .O(N__31454),
            .I(N__31297));
    Span4Mux_s1_h I__7382 (
            .O(N__31449),
            .I(N__31297));
    LocalMux I__7381 (
            .O(N__31440),
            .I(N__31292));
    LocalMux I__7380 (
            .O(N__31429),
            .I(N__31292));
    InMux I__7379 (
            .O(N__31428),
            .I(N__31281));
    InMux I__7378 (
            .O(N__31427),
            .I(N__31281));
    InMux I__7377 (
            .O(N__31426),
            .I(N__31281));
    InMux I__7376 (
            .O(N__31425),
            .I(N__31281));
    InMux I__7375 (
            .O(N__31424),
            .I(N__31281));
    Span4Mux_v I__7374 (
            .O(N__31421),
            .I(N__31274));
    LocalMux I__7373 (
            .O(N__31414),
            .I(N__31271));
    LocalMux I__7372 (
            .O(N__31409),
            .I(N__31264));
    LocalMux I__7371 (
            .O(N__31404),
            .I(N__31264));
    LocalMux I__7370 (
            .O(N__31399),
            .I(N__31264));
    InMux I__7369 (
            .O(N__31398),
            .I(N__31255));
    InMux I__7368 (
            .O(N__31395),
            .I(N__31255));
    InMux I__7367 (
            .O(N__31394),
            .I(N__31255));
    InMux I__7366 (
            .O(N__31393),
            .I(N__31255));
    InMux I__7365 (
            .O(N__31392),
            .I(N__31248));
    InMux I__7364 (
            .O(N__31391),
            .I(N__31248));
    InMux I__7363 (
            .O(N__31390),
            .I(N__31248));
    LocalMux I__7362 (
            .O(N__31387),
            .I(N__31245));
    InMux I__7361 (
            .O(N__31386),
            .I(N__31238));
    InMux I__7360 (
            .O(N__31385),
            .I(N__31238));
    InMux I__7359 (
            .O(N__31384),
            .I(N__31238));
    Span4Mux_s2_h I__7358 (
            .O(N__31381),
            .I(N__31231));
    Span4Mux_h I__7357 (
            .O(N__31378),
            .I(N__31231));
    LocalMux I__7356 (
            .O(N__31375),
            .I(N__31231));
    Span4Mux_v I__7355 (
            .O(N__31370),
            .I(N__31228));
    LocalMux I__7354 (
            .O(N__31359),
            .I(N__31225));
    InMux I__7353 (
            .O(N__31356),
            .I(N__31222));
    Span4Mux_h I__7352 (
            .O(N__31353),
            .I(N__31210));
    Span4Mux_h I__7351 (
            .O(N__31350),
            .I(N__31210));
    LocalMux I__7350 (
            .O(N__31343),
            .I(N__31210));
    InMux I__7349 (
            .O(N__31342),
            .I(N__31195));
    InMux I__7348 (
            .O(N__31341),
            .I(N__31195));
    InMux I__7347 (
            .O(N__31340),
            .I(N__31195));
    InMux I__7346 (
            .O(N__31339),
            .I(N__31195));
    InMux I__7345 (
            .O(N__31338),
            .I(N__31195));
    InMux I__7344 (
            .O(N__31337),
            .I(N__31195));
    InMux I__7343 (
            .O(N__31336),
            .I(N__31195));
    LocalMux I__7342 (
            .O(N__31327),
            .I(N__31192));
    InMux I__7341 (
            .O(N__31326),
            .I(N__31181));
    InMux I__7340 (
            .O(N__31325),
            .I(N__31181));
    InMux I__7339 (
            .O(N__31322),
            .I(N__31181));
    InMux I__7338 (
            .O(N__31321),
            .I(N__31181));
    InMux I__7337 (
            .O(N__31320),
            .I(N__31181));
    LocalMux I__7336 (
            .O(N__31317),
            .I(N__31176));
    Span4Mux_h I__7335 (
            .O(N__31306),
            .I(N__31176));
    CascadeMux I__7334 (
            .O(N__31305),
            .I(N__31169));
    Span4Mux_h I__7333 (
            .O(N__31302),
            .I(N__31166));
    Span4Mux_h I__7332 (
            .O(N__31297),
            .I(N__31159));
    Span4Mux_v I__7331 (
            .O(N__31292),
            .I(N__31159));
    LocalMux I__7330 (
            .O(N__31281),
            .I(N__31159));
    InMux I__7329 (
            .O(N__31280),
            .I(N__31150));
    InMux I__7328 (
            .O(N__31279),
            .I(N__31150));
    InMux I__7327 (
            .O(N__31278),
            .I(N__31150));
    InMux I__7326 (
            .O(N__31277),
            .I(N__31150));
    Span4Mux_h I__7325 (
            .O(N__31274),
            .I(N__31141));
    Span4Mux_v I__7324 (
            .O(N__31271),
            .I(N__31141));
    Span4Mux_v I__7323 (
            .O(N__31264),
            .I(N__31141));
    LocalMux I__7322 (
            .O(N__31255),
            .I(N__31141));
    LocalMux I__7321 (
            .O(N__31248),
            .I(N__31134));
    Span4Mux_v I__7320 (
            .O(N__31245),
            .I(N__31134));
    LocalMux I__7319 (
            .O(N__31238),
            .I(N__31134));
    Sp12to4 I__7318 (
            .O(N__31231),
            .I(N__31131));
    Span4Mux_h I__7317 (
            .O(N__31228),
            .I(N__31128));
    Span4Mux_h I__7316 (
            .O(N__31225),
            .I(N__31123));
    LocalMux I__7315 (
            .O(N__31222),
            .I(N__31123));
    InMux I__7314 (
            .O(N__31221),
            .I(N__31112));
    InMux I__7313 (
            .O(N__31220),
            .I(N__31112));
    InMux I__7312 (
            .O(N__31219),
            .I(N__31112));
    InMux I__7311 (
            .O(N__31218),
            .I(N__31112));
    InMux I__7310 (
            .O(N__31217),
            .I(N__31112));
    Span4Mux_v I__7309 (
            .O(N__31210),
            .I(N__31107));
    LocalMux I__7308 (
            .O(N__31195),
            .I(N__31107));
    Span4Mux_h I__7307 (
            .O(N__31192),
            .I(N__31100));
    LocalMux I__7306 (
            .O(N__31181),
            .I(N__31100));
    Span4Mux_v I__7305 (
            .O(N__31176),
            .I(N__31100));
    InMux I__7304 (
            .O(N__31175),
            .I(N__31089));
    InMux I__7303 (
            .O(N__31174),
            .I(N__31089));
    InMux I__7302 (
            .O(N__31173),
            .I(N__31089));
    InMux I__7301 (
            .O(N__31172),
            .I(N__31089));
    InMux I__7300 (
            .O(N__31169),
            .I(N__31089));
    Span4Mux_v I__7299 (
            .O(N__31166),
            .I(N__31078));
    Span4Mux_h I__7298 (
            .O(N__31159),
            .I(N__31078));
    LocalMux I__7297 (
            .O(N__31150),
            .I(N__31078));
    Span4Mux_h I__7296 (
            .O(N__31141),
            .I(N__31078));
    Span4Mux_h I__7295 (
            .O(N__31134),
            .I(N__31078));
    Odrv12 I__7294 (
            .O(N__31131),
            .I(instruction_9));
    Odrv4 I__7293 (
            .O(N__31128),
            .I(instruction_9));
    Odrv4 I__7292 (
            .O(N__31123),
            .I(instruction_9));
    LocalMux I__7291 (
            .O(N__31112),
            .I(instruction_9));
    Odrv4 I__7290 (
            .O(N__31107),
            .I(instruction_9));
    Odrv4 I__7289 (
            .O(N__31100),
            .I(instruction_9));
    LocalMux I__7288 (
            .O(N__31089),
            .I(instruction_9));
    Odrv4 I__7287 (
            .O(N__31078),
            .I(instruction_9));
    InMux I__7286 (
            .O(N__31061),
            .I(N__31057));
    InMux I__7285 (
            .O(N__31060),
            .I(N__31054));
    LocalMux I__7284 (
            .O(N__31057),
            .I(N__31049));
    LocalMux I__7283 (
            .O(N__31054),
            .I(N__31049));
    Span4Mux_v I__7282 (
            .O(N__31049),
            .I(N__31046));
    Odrv4 I__7281 (
            .O(N__31046),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_7 ));
    CascadeMux I__7280 (
            .O(N__31043),
            .I(N__31040));
    InMux I__7279 (
            .O(N__31040),
            .I(N__31036));
    InMux I__7278 (
            .O(N__31039),
            .I(N__31033));
    LocalMux I__7277 (
            .O(N__31036),
            .I(N__31028));
    LocalMux I__7276 (
            .O(N__31033),
            .I(N__31028));
    Span4Mux_v I__7275 (
            .O(N__31028),
            .I(N__31025));
    Odrv4 I__7274 (
            .O(N__31025),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_7 ));
    CascadeMux I__7273 (
            .O(N__31022),
            .I(N__31018));
    InMux I__7272 (
            .O(N__31021),
            .I(N__31010));
    InMux I__7271 (
            .O(N__31018),
            .I(N__31001));
    CascadeMux I__7270 (
            .O(N__31017),
            .I(N__30997));
    CascadeMux I__7269 (
            .O(N__31016),
            .I(N__30994));
    CascadeMux I__7268 (
            .O(N__31015),
            .I(N__30990));
    CascadeMux I__7267 (
            .O(N__31014),
            .I(N__30987));
    InMux I__7266 (
            .O(N__31013),
            .I(N__30976));
    LocalMux I__7265 (
            .O(N__31010),
            .I(N__30970));
    InMux I__7264 (
            .O(N__31009),
            .I(N__30967));
    InMux I__7263 (
            .O(N__31008),
            .I(N__30962));
    InMux I__7262 (
            .O(N__31007),
            .I(N__30962));
    InMux I__7261 (
            .O(N__31006),
            .I(N__30957));
    InMux I__7260 (
            .O(N__31005),
            .I(N__30957));
    InMux I__7259 (
            .O(N__31004),
            .I(N__30954));
    LocalMux I__7258 (
            .O(N__31001),
            .I(N__30951));
    InMux I__7257 (
            .O(N__31000),
            .I(N__30946));
    InMux I__7256 (
            .O(N__30997),
            .I(N__30946));
    InMux I__7255 (
            .O(N__30994),
            .I(N__30939));
    InMux I__7254 (
            .O(N__30993),
            .I(N__30936));
    InMux I__7253 (
            .O(N__30990),
            .I(N__30933));
    InMux I__7252 (
            .O(N__30987),
            .I(N__30928));
    InMux I__7251 (
            .O(N__30986),
            .I(N__30923));
    InMux I__7250 (
            .O(N__30985),
            .I(N__30923));
    InMux I__7249 (
            .O(N__30984),
            .I(N__30918));
    InMux I__7248 (
            .O(N__30983),
            .I(N__30911));
    InMux I__7247 (
            .O(N__30982),
            .I(N__30911));
    InMux I__7246 (
            .O(N__30981),
            .I(N__30904));
    InMux I__7245 (
            .O(N__30980),
            .I(N__30904));
    CascadeMux I__7244 (
            .O(N__30979),
            .I(N__30901));
    LocalMux I__7243 (
            .O(N__30976),
            .I(N__30895));
    InMux I__7242 (
            .O(N__30975),
            .I(N__30892));
    InMux I__7241 (
            .O(N__30974),
            .I(N__30887));
    InMux I__7240 (
            .O(N__30973),
            .I(N__30887));
    Span4Mux_s2_h I__7239 (
            .O(N__30970),
            .I(N__30882));
    LocalMux I__7238 (
            .O(N__30967),
            .I(N__30882));
    LocalMux I__7237 (
            .O(N__30962),
            .I(N__30877));
    LocalMux I__7236 (
            .O(N__30957),
            .I(N__30877));
    LocalMux I__7235 (
            .O(N__30954),
            .I(N__30870));
    Span4Mux_s3_v I__7234 (
            .O(N__30951),
            .I(N__30870));
    LocalMux I__7233 (
            .O(N__30946),
            .I(N__30870));
    InMux I__7232 (
            .O(N__30945),
            .I(N__30865));
    InMux I__7231 (
            .O(N__30944),
            .I(N__30865));
    CascadeMux I__7230 (
            .O(N__30943),
            .I(N__30861));
    CascadeMux I__7229 (
            .O(N__30942),
            .I(N__30856));
    LocalMux I__7228 (
            .O(N__30939),
            .I(N__30849));
    LocalMux I__7227 (
            .O(N__30936),
            .I(N__30849));
    LocalMux I__7226 (
            .O(N__30933),
            .I(N__30849));
    InMux I__7225 (
            .O(N__30932),
            .I(N__30838));
    InMux I__7224 (
            .O(N__30931),
            .I(N__30838));
    LocalMux I__7223 (
            .O(N__30928),
            .I(N__30830));
    LocalMux I__7222 (
            .O(N__30923),
            .I(N__30827));
    InMux I__7221 (
            .O(N__30922),
            .I(N__30824));
    CascadeMux I__7220 (
            .O(N__30921),
            .I(N__30819));
    LocalMux I__7219 (
            .O(N__30918),
            .I(N__30816));
    InMux I__7218 (
            .O(N__30917),
            .I(N__30813));
    InMux I__7217 (
            .O(N__30916),
            .I(N__30810));
    LocalMux I__7216 (
            .O(N__30911),
            .I(N__30807));
    InMux I__7215 (
            .O(N__30910),
            .I(N__30802));
    InMux I__7214 (
            .O(N__30909),
            .I(N__30802));
    LocalMux I__7213 (
            .O(N__30904),
            .I(N__30799));
    InMux I__7212 (
            .O(N__30901),
            .I(N__30794));
    InMux I__7211 (
            .O(N__30900),
            .I(N__30787));
    InMux I__7210 (
            .O(N__30899),
            .I(N__30787));
    InMux I__7209 (
            .O(N__30898),
            .I(N__30787));
    Span4Mux_s3_v I__7208 (
            .O(N__30895),
            .I(N__30780));
    LocalMux I__7207 (
            .O(N__30892),
            .I(N__30780));
    LocalMux I__7206 (
            .O(N__30887),
            .I(N__30780));
    Span4Mux_h I__7205 (
            .O(N__30882),
            .I(N__30771));
    Span4Mux_v I__7204 (
            .O(N__30877),
            .I(N__30771));
    Span4Mux_v I__7203 (
            .O(N__30870),
            .I(N__30771));
    LocalMux I__7202 (
            .O(N__30865),
            .I(N__30771));
    InMux I__7201 (
            .O(N__30864),
            .I(N__30768));
    InMux I__7200 (
            .O(N__30861),
            .I(N__30765));
    InMux I__7199 (
            .O(N__30860),
            .I(N__30760));
    InMux I__7198 (
            .O(N__30859),
            .I(N__30760));
    InMux I__7197 (
            .O(N__30856),
            .I(N__30757));
    Span4Mux_v I__7196 (
            .O(N__30849),
            .I(N__30754));
    InMux I__7195 (
            .O(N__30848),
            .I(N__30749));
    InMux I__7194 (
            .O(N__30847),
            .I(N__30749));
    InMux I__7193 (
            .O(N__30846),
            .I(N__30744));
    InMux I__7192 (
            .O(N__30845),
            .I(N__30744));
    CascadeMux I__7191 (
            .O(N__30844),
            .I(N__30741));
    CascadeMux I__7190 (
            .O(N__30843),
            .I(N__30738));
    LocalMux I__7189 (
            .O(N__30838),
            .I(N__30735));
    InMux I__7188 (
            .O(N__30837),
            .I(N__30730));
    InMux I__7187 (
            .O(N__30836),
            .I(N__30730));
    InMux I__7186 (
            .O(N__30835),
            .I(N__30723));
    InMux I__7185 (
            .O(N__30834),
            .I(N__30723));
    InMux I__7184 (
            .O(N__30833),
            .I(N__30723));
    Span4Mux_v I__7183 (
            .O(N__30830),
            .I(N__30716));
    Span4Mux_v I__7182 (
            .O(N__30827),
            .I(N__30716));
    LocalMux I__7181 (
            .O(N__30824),
            .I(N__30716));
    InMux I__7180 (
            .O(N__30823),
            .I(N__30709));
    InMux I__7179 (
            .O(N__30822),
            .I(N__30709));
    InMux I__7178 (
            .O(N__30819),
            .I(N__30709));
    Span4Mux_v I__7177 (
            .O(N__30816),
            .I(N__30704));
    LocalMux I__7176 (
            .O(N__30813),
            .I(N__30704));
    LocalMux I__7175 (
            .O(N__30810),
            .I(N__30699));
    Span4Mux_s3_v I__7174 (
            .O(N__30807),
            .I(N__30699));
    LocalMux I__7173 (
            .O(N__30802),
            .I(N__30694));
    Span4Mux_v I__7172 (
            .O(N__30799),
            .I(N__30694));
    InMux I__7171 (
            .O(N__30798),
            .I(N__30685));
    InMux I__7170 (
            .O(N__30797),
            .I(N__30685));
    LocalMux I__7169 (
            .O(N__30794),
            .I(N__30682));
    LocalMux I__7168 (
            .O(N__30787),
            .I(N__30675));
    Span4Mux_v I__7167 (
            .O(N__30780),
            .I(N__30675));
    Span4Mux_v I__7166 (
            .O(N__30771),
            .I(N__30675));
    LocalMux I__7165 (
            .O(N__30768),
            .I(N__30670));
    LocalMux I__7164 (
            .O(N__30765),
            .I(N__30670));
    LocalMux I__7163 (
            .O(N__30760),
            .I(N__30667));
    LocalMux I__7162 (
            .O(N__30757),
            .I(N__30660));
    Span4Mux_h I__7161 (
            .O(N__30754),
            .I(N__30660));
    LocalMux I__7160 (
            .O(N__30749),
            .I(N__30660));
    LocalMux I__7159 (
            .O(N__30744),
            .I(N__30653));
    InMux I__7158 (
            .O(N__30741),
            .I(N__30648));
    InMux I__7157 (
            .O(N__30738),
            .I(N__30648));
    Span4Mux_v I__7156 (
            .O(N__30735),
            .I(N__30637));
    LocalMux I__7155 (
            .O(N__30730),
            .I(N__30637));
    LocalMux I__7154 (
            .O(N__30723),
            .I(N__30637));
    Span4Mux_h I__7153 (
            .O(N__30716),
            .I(N__30637));
    LocalMux I__7152 (
            .O(N__30709),
            .I(N__30637));
    Span4Mux_h I__7151 (
            .O(N__30704),
            .I(N__30628));
    Span4Mux_v I__7150 (
            .O(N__30699),
            .I(N__30628));
    Span4Mux_v I__7149 (
            .O(N__30694),
            .I(N__30628));
    InMux I__7148 (
            .O(N__30693),
            .I(N__30623));
    InMux I__7147 (
            .O(N__30692),
            .I(N__30623));
    InMux I__7146 (
            .O(N__30691),
            .I(N__30618));
    InMux I__7145 (
            .O(N__30690),
            .I(N__30618));
    LocalMux I__7144 (
            .O(N__30685),
            .I(N__30609));
    Span4Mux_v I__7143 (
            .O(N__30682),
            .I(N__30609));
    Span4Mux_h I__7142 (
            .O(N__30675),
            .I(N__30609));
    Span4Mux_v I__7141 (
            .O(N__30670),
            .I(N__30609));
    Span4Mux_s2_h I__7140 (
            .O(N__30667),
            .I(N__30604));
    Span4Mux_h I__7139 (
            .O(N__30660),
            .I(N__30604));
    InMux I__7138 (
            .O(N__30659),
            .I(N__30595));
    InMux I__7137 (
            .O(N__30658),
            .I(N__30595));
    InMux I__7136 (
            .O(N__30657),
            .I(N__30595));
    InMux I__7135 (
            .O(N__30656),
            .I(N__30595));
    Span4Mux_v I__7134 (
            .O(N__30653),
            .I(N__30588));
    LocalMux I__7133 (
            .O(N__30648),
            .I(N__30588));
    Span4Mux_h I__7132 (
            .O(N__30637),
            .I(N__30588));
    InMux I__7131 (
            .O(N__30636),
            .I(N__30583));
    InMux I__7130 (
            .O(N__30635),
            .I(N__30583));
    Odrv4 I__7129 (
            .O(N__30628),
            .I(instruction_8));
    LocalMux I__7128 (
            .O(N__30623),
            .I(instruction_8));
    LocalMux I__7127 (
            .O(N__30618),
            .I(instruction_8));
    Odrv4 I__7126 (
            .O(N__30609),
            .I(instruction_8));
    Odrv4 I__7125 (
            .O(N__30604),
            .I(instruction_8));
    LocalMux I__7124 (
            .O(N__30595),
            .I(instruction_8));
    Odrv4 I__7123 (
            .O(N__30588),
            .I(instruction_8));
    LocalMux I__7122 (
            .O(N__30583),
            .I(instruction_8));
    InMux I__7121 (
            .O(N__30566),
            .I(N__30563));
    LocalMux I__7120 (
            .O(N__30563),
            .I(N__30560));
    Odrv12 I__7119 (
            .O(N__30560),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_7 ));
    InMux I__7118 (
            .O(N__30557),
            .I(N__30554));
    LocalMux I__7117 (
            .O(N__30554),
            .I(N__30550));
    InMux I__7116 (
            .O(N__30553),
            .I(N__30547));
    Span4Mux_v I__7115 (
            .O(N__30550),
            .I(N__30544));
    LocalMux I__7114 (
            .O(N__30547),
            .I(N__30541));
    Odrv4 I__7113 (
            .O(N__30544),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0 ));
    Odrv12 I__7112 (
            .O(N__30541),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0 ));
    InMux I__7111 (
            .O(N__30536),
            .I(N__30532));
    InMux I__7110 (
            .O(N__30535),
            .I(N__30529));
    LocalMux I__7109 (
            .O(N__30532),
            .I(N__30524));
    LocalMux I__7108 (
            .O(N__30529),
            .I(N__30524));
    Span4Mux_v I__7107 (
            .O(N__30524),
            .I(N__30521));
    Odrv4 I__7106 (
            .O(N__30521),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_3 ));
    CascadeMux I__7105 (
            .O(N__30518),
            .I(N__30515));
    InMux I__7104 (
            .O(N__30515),
            .I(N__30511));
    CascadeMux I__7103 (
            .O(N__30514),
            .I(N__30504));
    LocalMux I__7102 (
            .O(N__30511),
            .I(N__30501));
    CascadeMux I__7101 (
            .O(N__30510),
            .I(N__30495));
    CascadeMux I__7100 (
            .O(N__30509),
            .I(N__30486));
    CascadeMux I__7099 (
            .O(N__30508),
            .I(N__30482));
    CascadeMux I__7098 (
            .O(N__30507),
            .I(N__30478));
    InMux I__7097 (
            .O(N__30504),
            .I(N__30474));
    Span4Mux_s2_h I__7096 (
            .O(N__30501),
            .I(N__30468));
    InMux I__7095 (
            .O(N__30500),
            .I(N__30465));
    CascadeMux I__7094 (
            .O(N__30499),
            .I(N__30458));
    CascadeMux I__7093 (
            .O(N__30498),
            .I(N__30455));
    InMux I__7092 (
            .O(N__30495),
            .I(N__30452));
    InMux I__7091 (
            .O(N__30494),
            .I(N__30449));
    InMux I__7090 (
            .O(N__30493),
            .I(N__30445));
    CascadeMux I__7089 (
            .O(N__30492),
            .I(N__30441));
    CascadeMux I__7088 (
            .O(N__30491),
            .I(N__30436));
    CascadeMux I__7087 (
            .O(N__30490),
            .I(N__30433));
    InMux I__7086 (
            .O(N__30489),
            .I(N__30430));
    InMux I__7085 (
            .O(N__30486),
            .I(N__30427));
    InMux I__7084 (
            .O(N__30485),
            .I(N__30424));
    InMux I__7083 (
            .O(N__30482),
            .I(N__30421));
    InMux I__7082 (
            .O(N__30481),
            .I(N__30418));
    InMux I__7081 (
            .O(N__30478),
            .I(N__30415));
    InMux I__7080 (
            .O(N__30477),
            .I(N__30412));
    LocalMux I__7079 (
            .O(N__30474),
            .I(N__30409));
    CascadeMux I__7078 (
            .O(N__30473),
            .I(N__30406));
    CascadeMux I__7077 (
            .O(N__30472),
            .I(N__30403));
    CascadeMux I__7076 (
            .O(N__30471),
            .I(N__30400));
    Span4Mux_v I__7075 (
            .O(N__30468),
            .I(N__30395));
    LocalMux I__7074 (
            .O(N__30465),
            .I(N__30395));
    InMux I__7073 (
            .O(N__30464),
            .I(N__30391));
    CascadeMux I__7072 (
            .O(N__30463),
            .I(N__30387));
    CascadeMux I__7071 (
            .O(N__30462),
            .I(N__30383));
    InMux I__7070 (
            .O(N__30461),
            .I(N__30380));
    InMux I__7069 (
            .O(N__30458),
            .I(N__30377));
    InMux I__7068 (
            .O(N__30455),
            .I(N__30374));
    LocalMux I__7067 (
            .O(N__30452),
            .I(N__30371));
    LocalMux I__7066 (
            .O(N__30449),
            .I(N__30368));
    InMux I__7065 (
            .O(N__30448),
            .I(N__30365));
    LocalMux I__7064 (
            .O(N__30445),
            .I(N__30362));
    CascadeMux I__7063 (
            .O(N__30444),
            .I(N__30359));
    InMux I__7062 (
            .O(N__30441),
            .I(N__30356));
    InMux I__7061 (
            .O(N__30440),
            .I(N__30353));
    InMux I__7060 (
            .O(N__30439),
            .I(N__30350));
    InMux I__7059 (
            .O(N__30436),
            .I(N__30347));
    InMux I__7058 (
            .O(N__30433),
            .I(N__30344));
    LocalMux I__7057 (
            .O(N__30430),
            .I(N__30341));
    LocalMux I__7056 (
            .O(N__30427),
            .I(N__30338));
    LocalMux I__7055 (
            .O(N__30424),
            .I(N__30335));
    LocalMux I__7054 (
            .O(N__30421),
            .I(N__30332));
    LocalMux I__7053 (
            .O(N__30418),
            .I(N__30323));
    LocalMux I__7052 (
            .O(N__30415),
            .I(N__30323));
    LocalMux I__7051 (
            .O(N__30412),
            .I(N__30323));
    Span4Mux_v I__7050 (
            .O(N__30409),
            .I(N__30323));
    InMux I__7049 (
            .O(N__30406),
            .I(N__30320));
    InMux I__7048 (
            .O(N__30403),
            .I(N__30317));
    InMux I__7047 (
            .O(N__30400),
            .I(N__30314));
    Span4Mux_h I__7046 (
            .O(N__30395),
            .I(N__30311));
    InMux I__7045 (
            .O(N__30394),
            .I(N__30308));
    LocalMux I__7044 (
            .O(N__30391),
            .I(N__30305));
    InMux I__7043 (
            .O(N__30390),
            .I(N__30302));
    InMux I__7042 (
            .O(N__30387),
            .I(N__30299));
    InMux I__7041 (
            .O(N__30386),
            .I(N__30296));
    InMux I__7040 (
            .O(N__30383),
            .I(N__30293));
    LocalMux I__7039 (
            .O(N__30380),
            .I(N__30288));
    LocalMux I__7038 (
            .O(N__30377),
            .I(N__30288));
    LocalMux I__7037 (
            .O(N__30374),
            .I(N__30281));
    Span4Mux_v I__7036 (
            .O(N__30371),
            .I(N__30281));
    Span4Mux_v I__7035 (
            .O(N__30368),
            .I(N__30281));
    LocalMux I__7034 (
            .O(N__30365),
            .I(N__30276));
    Span4Mux_s3_v I__7033 (
            .O(N__30362),
            .I(N__30276));
    InMux I__7032 (
            .O(N__30359),
            .I(N__30273));
    LocalMux I__7031 (
            .O(N__30356),
            .I(N__30270));
    LocalMux I__7030 (
            .O(N__30353),
            .I(N__30254));
    LocalMux I__7029 (
            .O(N__30350),
            .I(N__30254));
    LocalMux I__7028 (
            .O(N__30347),
            .I(N__30254));
    LocalMux I__7027 (
            .O(N__30344),
            .I(N__30254));
    Span4Mux_v I__7026 (
            .O(N__30341),
            .I(N__30254));
    Span4Mux_h I__7025 (
            .O(N__30338),
            .I(N__30254));
    Span4Mux_s2_v I__7024 (
            .O(N__30335),
            .I(N__30254));
    Span4Mux_s3_h I__7023 (
            .O(N__30332),
            .I(N__30251));
    Span4Mux_v I__7022 (
            .O(N__30323),
            .I(N__30248));
    LocalMux I__7021 (
            .O(N__30320),
            .I(N__30241));
    LocalMux I__7020 (
            .O(N__30317),
            .I(N__30241));
    LocalMux I__7019 (
            .O(N__30314),
            .I(N__30241));
    Sp12to4 I__7018 (
            .O(N__30311),
            .I(N__30238));
    LocalMux I__7017 (
            .O(N__30308),
            .I(N__30235));
    Span4Mux_s2_v I__7016 (
            .O(N__30305),
            .I(N__30232));
    LocalMux I__7015 (
            .O(N__30302),
            .I(N__30229));
    LocalMux I__7014 (
            .O(N__30299),
            .I(N__30224));
    LocalMux I__7013 (
            .O(N__30296),
            .I(N__30224));
    LocalMux I__7012 (
            .O(N__30293),
            .I(N__30219));
    Span4Mux_v I__7011 (
            .O(N__30288),
            .I(N__30219));
    Span4Mux_v I__7010 (
            .O(N__30281),
            .I(N__30214));
    Span4Mux_v I__7009 (
            .O(N__30276),
            .I(N__30214));
    LocalMux I__7008 (
            .O(N__30273),
            .I(N__30211));
    Span4Mux_s2_h I__7007 (
            .O(N__30270),
            .I(N__30208));
    InMux I__7006 (
            .O(N__30269),
            .I(N__30204));
    Span4Mux_v I__7005 (
            .O(N__30254),
            .I(N__30197));
    Span4Mux_v I__7004 (
            .O(N__30251),
            .I(N__30197));
    Span4Mux_h I__7003 (
            .O(N__30248),
            .I(N__30197));
    Span12Mux_s6_h I__7002 (
            .O(N__30241),
            .I(N__30192));
    Span12Mux_s3_v I__7001 (
            .O(N__30238),
            .I(N__30192));
    Span4Mux_h I__7000 (
            .O(N__30235),
            .I(N__30187));
    Span4Mux_v I__6999 (
            .O(N__30232),
            .I(N__30187));
    Span4Mux_v I__6998 (
            .O(N__30229),
            .I(N__30178));
    Span4Mux_v I__6997 (
            .O(N__30224),
            .I(N__30178));
    Span4Mux_h I__6996 (
            .O(N__30219),
            .I(N__30178));
    Span4Mux_h I__6995 (
            .O(N__30214),
            .I(N__30178));
    Span4Mux_v I__6994 (
            .O(N__30211),
            .I(N__30173));
    Span4Mux_v I__6993 (
            .O(N__30208),
            .I(N__30173));
    InMux I__6992 (
            .O(N__30207),
            .I(N__30170));
    LocalMux I__6991 (
            .O(N__30204),
            .I(\processor_zipi8.arith_logical_result_5 ));
    Odrv4 I__6990 (
            .O(N__30197),
            .I(\processor_zipi8.arith_logical_result_5 ));
    Odrv12 I__6989 (
            .O(N__30192),
            .I(\processor_zipi8.arith_logical_result_5 ));
    Odrv4 I__6988 (
            .O(N__30187),
            .I(\processor_zipi8.arith_logical_result_5 ));
    Odrv4 I__6987 (
            .O(N__30178),
            .I(\processor_zipi8.arith_logical_result_5 ));
    Odrv4 I__6986 (
            .O(N__30173),
            .I(\processor_zipi8.arith_logical_result_5 ));
    LocalMux I__6985 (
            .O(N__30170),
            .I(\processor_zipi8.arith_logical_result_5 ));
    CascadeMux I__6984 (
            .O(N__30155),
            .I(N__30151));
    InMux I__6983 (
            .O(N__30154),
            .I(N__30141));
    InMux I__6982 (
            .O(N__30151),
            .I(N__30138));
    CascadeMux I__6981 (
            .O(N__30150),
            .I(N__30131));
    InMux I__6980 (
            .O(N__30149),
            .I(N__30128));
    InMux I__6979 (
            .O(N__30148),
            .I(N__30125));
    InMux I__6978 (
            .O(N__30147),
            .I(N__30122));
    CascadeMux I__6977 (
            .O(N__30146),
            .I(N__30118));
    InMux I__6976 (
            .O(N__30145),
            .I(N__30112));
    InMux I__6975 (
            .O(N__30144),
            .I(N__30109));
    LocalMux I__6974 (
            .O(N__30141),
            .I(N__30106));
    LocalMux I__6973 (
            .O(N__30138),
            .I(N__30103));
    CascadeMux I__6972 (
            .O(N__30137),
            .I(N__30100));
    CascadeMux I__6971 (
            .O(N__30136),
            .I(N__30097));
    CascadeMux I__6970 (
            .O(N__30135),
            .I(N__30094));
    CascadeMux I__6969 (
            .O(N__30134),
            .I(N__30091));
    InMux I__6968 (
            .O(N__30131),
            .I(N__30085));
    LocalMux I__6967 (
            .O(N__30128),
            .I(N__30082));
    LocalMux I__6966 (
            .O(N__30125),
            .I(N__30077));
    LocalMux I__6965 (
            .O(N__30122),
            .I(N__30077));
    CascadeMux I__6964 (
            .O(N__30121),
            .I(N__30073));
    InMux I__6963 (
            .O(N__30118),
            .I(N__30070));
    InMux I__6962 (
            .O(N__30117),
            .I(N__30064));
    InMux I__6961 (
            .O(N__30116),
            .I(N__30061));
    InMux I__6960 (
            .O(N__30115),
            .I(N__30058));
    LocalMux I__6959 (
            .O(N__30112),
            .I(N__30048));
    LocalMux I__6958 (
            .O(N__30109),
            .I(N__30048));
    Span4Mux_s2_h I__6957 (
            .O(N__30106),
            .I(N__30048));
    Span4Mux_s3_v I__6956 (
            .O(N__30103),
            .I(N__30048));
    InMux I__6955 (
            .O(N__30100),
            .I(N__30045));
    InMux I__6954 (
            .O(N__30097),
            .I(N__30041));
    InMux I__6953 (
            .O(N__30094),
            .I(N__30038));
    InMux I__6952 (
            .O(N__30091),
            .I(N__30035));
    CascadeMux I__6951 (
            .O(N__30090),
            .I(N__30031));
    InMux I__6950 (
            .O(N__30089),
            .I(N__30028));
    CascadeMux I__6949 (
            .O(N__30088),
            .I(N__30025));
    LocalMux I__6948 (
            .O(N__30085),
            .I(N__30021));
    Span4Mux_v I__6947 (
            .O(N__30082),
            .I(N__30016));
    Span4Mux_v I__6946 (
            .O(N__30077),
            .I(N__30016));
    InMux I__6945 (
            .O(N__30076),
            .I(N__30013));
    InMux I__6944 (
            .O(N__30073),
            .I(N__30010));
    LocalMux I__6943 (
            .O(N__30070),
            .I(N__30007));
    InMux I__6942 (
            .O(N__30069),
            .I(N__30004));
    InMux I__6941 (
            .O(N__30068),
            .I(N__30001));
    InMux I__6940 (
            .O(N__30067),
            .I(N__29998));
    LocalMux I__6939 (
            .O(N__30064),
            .I(N__29993));
    LocalMux I__6938 (
            .O(N__30061),
            .I(N__29993));
    LocalMux I__6937 (
            .O(N__30058),
            .I(N__29990));
    InMux I__6936 (
            .O(N__30057),
            .I(N__29987));
    Span4Mux_h I__6935 (
            .O(N__30048),
            .I(N__29982));
    LocalMux I__6934 (
            .O(N__30045),
            .I(N__29982));
    CascadeMux I__6933 (
            .O(N__30044),
            .I(N__29979));
    LocalMux I__6932 (
            .O(N__30041),
            .I(N__29974));
    LocalMux I__6931 (
            .O(N__30038),
            .I(N__29974));
    LocalMux I__6930 (
            .O(N__30035),
            .I(N__29971));
    InMux I__6929 (
            .O(N__30034),
            .I(N__29968));
    InMux I__6928 (
            .O(N__30031),
            .I(N__29965));
    LocalMux I__6927 (
            .O(N__30028),
            .I(N__29962));
    InMux I__6926 (
            .O(N__30025),
            .I(N__29959));
    InMux I__6925 (
            .O(N__30024),
            .I(N__29956));
    Span4Mux_v I__6924 (
            .O(N__30021),
            .I(N__29953));
    Span4Mux_s0_h I__6923 (
            .O(N__30016),
            .I(N__29947));
    LocalMux I__6922 (
            .O(N__30013),
            .I(N__29944));
    LocalMux I__6921 (
            .O(N__30010),
            .I(N__29937));
    Span4Mux_s3_v I__6920 (
            .O(N__30007),
            .I(N__29937));
    LocalMux I__6919 (
            .O(N__30004),
            .I(N__29937));
    LocalMux I__6918 (
            .O(N__30001),
            .I(N__29928));
    LocalMux I__6917 (
            .O(N__29998),
            .I(N__29928));
    Span4Mux_v I__6916 (
            .O(N__29993),
            .I(N__29928));
    Span4Mux_v I__6915 (
            .O(N__29990),
            .I(N__29928));
    LocalMux I__6914 (
            .O(N__29987),
            .I(N__29923));
    Span4Mux_v I__6913 (
            .O(N__29982),
            .I(N__29923));
    InMux I__6912 (
            .O(N__29979),
            .I(N__29920));
    Span4Mux_s1_h I__6911 (
            .O(N__29974),
            .I(N__29917));
    Span4Mux_s2_v I__6910 (
            .O(N__29971),
            .I(N__29914));
    LocalMux I__6909 (
            .O(N__29968),
            .I(N__29911));
    LocalMux I__6908 (
            .O(N__29965),
            .I(N__29908));
    Span4Mux_h I__6907 (
            .O(N__29962),
            .I(N__29901));
    LocalMux I__6906 (
            .O(N__29959),
            .I(N__29901));
    LocalMux I__6905 (
            .O(N__29956),
            .I(N__29901));
    Span4Mux_h I__6904 (
            .O(N__29953),
            .I(N__29898));
    InMux I__6903 (
            .O(N__29952),
            .I(N__29895));
    InMux I__6902 (
            .O(N__29951),
            .I(N__29891));
    InMux I__6901 (
            .O(N__29950),
            .I(N__29888));
    Span4Mux_h I__6900 (
            .O(N__29947),
            .I(N__29885));
    Span4Mux_v I__6899 (
            .O(N__29944),
            .I(N__29878));
    Span4Mux_v I__6898 (
            .O(N__29937),
            .I(N__29878));
    Span4Mux_v I__6897 (
            .O(N__29928),
            .I(N__29878));
    Span4Mux_h I__6896 (
            .O(N__29923),
            .I(N__29875));
    LocalMux I__6895 (
            .O(N__29920),
            .I(N__29866));
    Span4Mux_h I__6894 (
            .O(N__29917),
            .I(N__29866));
    Span4Mux_v I__6893 (
            .O(N__29914),
            .I(N__29866));
    Span4Mux_v I__6892 (
            .O(N__29911),
            .I(N__29866));
    Span4Mux_h I__6891 (
            .O(N__29908),
            .I(N__29861));
    Span4Mux_v I__6890 (
            .O(N__29901),
            .I(N__29861));
    Span4Mux_h I__6889 (
            .O(N__29898),
            .I(N__29856));
    LocalMux I__6888 (
            .O(N__29895),
            .I(N__29856));
    InMux I__6887 (
            .O(N__29894),
            .I(N__29853));
    LocalMux I__6886 (
            .O(N__29891),
            .I(N__29848));
    LocalMux I__6885 (
            .O(N__29888),
            .I(N__29848));
    Span4Mux_h I__6884 (
            .O(N__29885),
            .I(N__29845));
    Sp12to4 I__6883 (
            .O(N__29878),
            .I(N__29842));
    Span4Mux_s1_h I__6882 (
            .O(N__29875),
            .I(N__29839));
    Span4Mux_h I__6881 (
            .O(N__29866),
            .I(N__29834));
    Span4Mux_h I__6880 (
            .O(N__29861),
            .I(N__29834));
    Span4Mux_v I__6879 (
            .O(N__29856),
            .I(N__29831));
    LocalMux I__6878 (
            .O(N__29853),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ));
    Odrv4 I__6877 (
            .O(N__29848),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ));
    Odrv4 I__6876 (
            .O(N__29845),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ));
    Odrv12 I__6875 (
            .O(N__29842),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ));
    Odrv4 I__6874 (
            .O(N__29839),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ));
    Odrv4 I__6873 (
            .O(N__29834),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ));
    Odrv4 I__6872 (
            .O(N__29831),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ));
    CascadeMux I__6871 (
            .O(N__29816),
            .I(N__29813));
    InMux I__6870 (
            .O(N__29813),
            .I(N__29809));
    InMux I__6869 (
            .O(N__29812),
            .I(N__29806));
    LocalMux I__6868 (
            .O(N__29809),
            .I(N__29803));
    LocalMux I__6867 (
            .O(N__29806),
            .I(N__29800));
    Span4Mux_v I__6866 (
            .O(N__29803),
            .I(N__29797));
    Span4Mux_v I__6865 (
            .O(N__29800),
            .I(N__29794));
    Span4Mux_h I__6864 (
            .O(N__29797),
            .I(N__29791));
    Sp12to4 I__6863 (
            .O(N__29794),
            .I(N__29788));
    Odrv4 I__6862 (
            .O(N__29791),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5 ));
    Odrv12 I__6861 (
            .O(N__29788),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5 ));
    CascadeMux I__6860 (
            .O(N__29783),
            .I(N__29777));
    CascadeMux I__6859 (
            .O(N__29782),
            .I(N__29774));
    InMux I__6858 (
            .O(N__29781),
            .I(N__29765));
    CascadeMux I__6857 (
            .O(N__29780),
            .I(N__29761));
    InMux I__6856 (
            .O(N__29777),
            .I(N__29758));
    InMux I__6855 (
            .O(N__29774),
            .I(N__29755));
    CascadeMux I__6854 (
            .O(N__29773),
            .I(N__29752));
    InMux I__6853 (
            .O(N__29772),
            .I(N__29748));
    InMux I__6852 (
            .O(N__29771),
            .I(N__29745));
    CascadeMux I__6851 (
            .O(N__29770),
            .I(N__29740));
    CascadeMux I__6850 (
            .O(N__29769),
            .I(N__29737));
    CascadeMux I__6849 (
            .O(N__29768),
            .I(N__29732));
    LocalMux I__6848 (
            .O(N__29765),
            .I(N__29729));
    InMux I__6847 (
            .O(N__29764),
            .I(N__29726));
    InMux I__6846 (
            .O(N__29761),
            .I(N__29723));
    LocalMux I__6845 (
            .O(N__29758),
            .I(N__29717));
    LocalMux I__6844 (
            .O(N__29755),
            .I(N__29717));
    InMux I__6843 (
            .O(N__29752),
            .I(N__29714));
    InMux I__6842 (
            .O(N__29751),
            .I(N__29711));
    LocalMux I__6841 (
            .O(N__29748),
            .I(N__29701));
    LocalMux I__6840 (
            .O(N__29745),
            .I(N__29698));
    InMux I__6839 (
            .O(N__29744),
            .I(N__29695));
    InMux I__6838 (
            .O(N__29743),
            .I(N__29692));
    InMux I__6837 (
            .O(N__29740),
            .I(N__29688));
    InMux I__6836 (
            .O(N__29737),
            .I(N__29685));
    CascadeMux I__6835 (
            .O(N__29736),
            .I(N__29681));
    InMux I__6834 (
            .O(N__29735),
            .I(N__29678));
    InMux I__6833 (
            .O(N__29732),
            .I(N__29672));
    Span4Mux_s3_v I__6832 (
            .O(N__29729),
            .I(N__29665));
    LocalMux I__6831 (
            .O(N__29726),
            .I(N__29665));
    LocalMux I__6830 (
            .O(N__29723),
            .I(N__29665));
    InMux I__6829 (
            .O(N__29722),
            .I(N__29662));
    Span4Mux_v I__6828 (
            .O(N__29717),
            .I(N__29659));
    LocalMux I__6827 (
            .O(N__29714),
            .I(N__29656));
    LocalMux I__6826 (
            .O(N__29711),
            .I(N__29653));
    InMux I__6825 (
            .O(N__29710),
            .I(N__29650));
    InMux I__6824 (
            .O(N__29709),
            .I(N__29647));
    InMux I__6823 (
            .O(N__29708),
            .I(N__29644));
    InMux I__6822 (
            .O(N__29707),
            .I(N__29639));
    InMux I__6821 (
            .O(N__29706),
            .I(N__29636));
    CascadeMux I__6820 (
            .O(N__29705),
            .I(N__29633));
    CascadeMux I__6819 (
            .O(N__29704),
            .I(N__29630));
    Span4Mux_s2_h I__6818 (
            .O(N__29701),
            .I(N__29621));
    Span4Mux_s3_v I__6817 (
            .O(N__29698),
            .I(N__29621));
    LocalMux I__6816 (
            .O(N__29695),
            .I(N__29621));
    LocalMux I__6815 (
            .O(N__29692),
            .I(N__29621));
    InMux I__6814 (
            .O(N__29691),
            .I(N__29618));
    LocalMux I__6813 (
            .O(N__29688),
            .I(N__29615));
    LocalMux I__6812 (
            .O(N__29685),
            .I(N__29612));
    InMux I__6811 (
            .O(N__29684),
            .I(N__29609));
    InMux I__6810 (
            .O(N__29681),
            .I(N__29606));
    LocalMux I__6809 (
            .O(N__29678),
            .I(N__29603));
    InMux I__6808 (
            .O(N__29677),
            .I(N__29600));
    InMux I__6807 (
            .O(N__29676),
            .I(N__29597));
    InMux I__6806 (
            .O(N__29675),
            .I(N__29594));
    LocalMux I__6805 (
            .O(N__29672),
            .I(N__29591));
    Span4Mux_v I__6804 (
            .O(N__29665),
            .I(N__29586));
    LocalMux I__6803 (
            .O(N__29662),
            .I(N__29586));
    Span4Mux_v I__6802 (
            .O(N__29659),
            .I(N__29581));
    Span4Mux_s3_v I__6801 (
            .O(N__29656),
            .I(N__29581));
    Span4Mux_s0_h I__6800 (
            .O(N__29653),
            .I(N__29572));
    LocalMux I__6799 (
            .O(N__29650),
            .I(N__29572));
    LocalMux I__6798 (
            .O(N__29647),
            .I(N__29572));
    LocalMux I__6797 (
            .O(N__29644),
            .I(N__29572));
    CascadeMux I__6796 (
            .O(N__29643),
            .I(N__29569));
    InMux I__6795 (
            .O(N__29642),
            .I(N__29566));
    LocalMux I__6794 (
            .O(N__29639),
            .I(N__29561));
    LocalMux I__6793 (
            .O(N__29636),
            .I(N__29561));
    InMux I__6792 (
            .O(N__29633),
            .I(N__29558));
    InMux I__6791 (
            .O(N__29630),
            .I(N__29555));
    Span4Mux_h I__6790 (
            .O(N__29621),
            .I(N__29548));
    LocalMux I__6789 (
            .O(N__29618),
            .I(N__29548));
    Span4Mux_v I__6788 (
            .O(N__29615),
            .I(N__29541));
    Span4Mux_v I__6787 (
            .O(N__29612),
            .I(N__29541));
    LocalMux I__6786 (
            .O(N__29609),
            .I(N__29541));
    LocalMux I__6785 (
            .O(N__29606),
            .I(N__29538));
    Span4Mux_h I__6784 (
            .O(N__29603),
            .I(N__29529));
    LocalMux I__6783 (
            .O(N__29600),
            .I(N__29529));
    LocalMux I__6782 (
            .O(N__29597),
            .I(N__29529));
    LocalMux I__6781 (
            .O(N__29594),
            .I(N__29529));
    Span4Mux_s3_h I__6780 (
            .O(N__29591),
            .I(N__29524));
    Span4Mux_v I__6779 (
            .O(N__29586),
            .I(N__29524));
    Span4Mux_v I__6778 (
            .O(N__29581),
            .I(N__29519));
    Span4Mux_v I__6777 (
            .O(N__29572),
            .I(N__29519));
    InMux I__6776 (
            .O(N__29569),
            .I(N__29516));
    LocalMux I__6775 (
            .O(N__29566),
            .I(N__29513));
    Span4Mux_v I__6774 (
            .O(N__29561),
            .I(N__29506));
    LocalMux I__6773 (
            .O(N__29558),
            .I(N__29506));
    LocalMux I__6772 (
            .O(N__29555),
            .I(N__29506));
    InMux I__6771 (
            .O(N__29554),
            .I(N__29503));
    InMux I__6770 (
            .O(N__29553),
            .I(N__29500));
    Span4Mux_h I__6769 (
            .O(N__29548),
            .I(N__29496));
    Span4Mux_h I__6768 (
            .O(N__29541),
            .I(N__29493));
    Span4Mux_v I__6767 (
            .O(N__29538),
            .I(N__29490));
    Span4Mux_v I__6766 (
            .O(N__29529),
            .I(N__29485));
    Span4Mux_h I__6765 (
            .O(N__29524),
            .I(N__29485));
    Sp12to4 I__6764 (
            .O(N__29519),
            .I(N__29480));
    LocalMux I__6763 (
            .O(N__29516),
            .I(N__29480));
    Span4Mux_h I__6762 (
            .O(N__29513),
            .I(N__29477));
    Span4Mux_h I__6761 (
            .O(N__29506),
            .I(N__29470));
    LocalMux I__6760 (
            .O(N__29503),
            .I(N__29470));
    LocalMux I__6759 (
            .O(N__29500),
            .I(N__29470));
    InMux I__6758 (
            .O(N__29499),
            .I(N__29467));
    Span4Mux_v I__6757 (
            .O(N__29496),
            .I(N__29460));
    Span4Mux_h I__6756 (
            .O(N__29493),
            .I(N__29460));
    Span4Mux_h I__6755 (
            .O(N__29490),
            .I(N__29460));
    Odrv4 I__6754 (
            .O(N__29485),
            .I(\processor_zipi8.arith_logical_result_6 ));
    Odrv12 I__6753 (
            .O(N__29480),
            .I(\processor_zipi8.arith_logical_result_6 ));
    Odrv4 I__6752 (
            .O(N__29477),
            .I(\processor_zipi8.arith_logical_result_6 ));
    Odrv4 I__6751 (
            .O(N__29470),
            .I(\processor_zipi8.arith_logical_result_6 ));
    LocalMux I__6750 (
            .O(N__29467),
            .I(\processor_zipi8.arith_logical_result_6 ));
    Odrv4 I__6749 (
            .O(N__29460),
            .I(\processor_zipi8.arith_logical_result_6 ));
    InMux I__6748 (
            .O(N__29447),
            .I(N__29442));
    CascadeMux I__6747 (
            .O(N__29446),
            .I(N__29439));
    InMux I__6746 (
            .O(N__29445),
            .I(N__29434));
    LocalMux I__6745 (
            .O(N__29442),
            .I(N__29431));
    InMux I__6744 (
            .O(N__29439),
            .I(N__29428));
    InMux I__6743 (
            .O(N__29438),
            .I(N__29425));
    CascadeMux I__6742 (
            .O(N__29437),
            .I(N__29422));
    LocalMux I__6741 (
            .O(N__29434),
            .I(N__29415));
    Span4Mux_s1_v I__6740 (
            .O(N__29431),
            .I(N__29415));
    LocalMux I__6739 (
            .O(N__29428),
            .I(N__29415));
    LocalMux I__6738 (
            .O(N__29425),
            .I(N__29412));
    InMux I__6737 (
            .O(N__29422),
            .I(N__29409));
    Span4Mux_h I__6736 (
            .O(N__29415),
            .I(N__29399));
    Span4Mux_v I__6735 (
            .O(N__29412),
            .I(N__29399));
    LocalMux I__6734 (
            .O(N__29409),
            .I(N__29399));
    CascadeMux I__6733 (
            .O(N__29408),
            .I(N__29390));
    CascadeMux I__6732 (
            .O(N__29407),
            .I(N__29387));
    CascadeMux I__6731 (
            .O(N__29406),
            .I(N__29384));
    Span4Mux_v I__6730 (
            .O(N__29399),
            .I(N__29381));
    InMux I__6729 (
            .O(N__29398),
            .I(N__29378));
    CascadeMux I__6728 (
            .O(N__29397),
            .I(N__29375));
    InMux I__6727 (
            .O(N__29396),
            .I(N__29372));
    CascadeMux I__6726 (
            .O(N__29395),
            .I(N__29361));
    CascadeMux I__6725 (
            .O(N__29394),
            .I(N__29358));
    InMux I__6724 (
            .O(N__29393),
            .I(N__29353));
    InMux I__6723 (
            .O(N__29390),
            .I(N__29350));
    InMux I__6722 (
            .O(N__29387),
            .I(N__29347));
    InMux I__6721 (
            .O(N__29384),
            .I(N__29344));
    Span4Mux_s0_h I__6720 (
            .O(N__29381),
            .I(N__29339));
    LocalMux I__6719 (
            .O(N__29378),
            .I(N__29339));
    InMux I__6718 (
            .O(N__29375),
            .I(N__29336));
    LocalMux I__6717 (
            .O(N__29372),
            .I(N__29333));
    InMux I__6716 (
            .O(N__29371),
            .I(N__29330));
    CascadeMux I__6715 (
            .O(N__29370),
            .I(N__29326));
    CascadeMux I__6714 (
            .O(N__29369),
            .I(N__29323));
    CascadeMux I__6713 (
            .O(N__29368),
            .I(N__29320));
    CascadeMux I__6712 (
            .O(N__29367),
            .I(N__29317));
    CascadeMux I__6711 (
            .O(N__29366),
            .I(N__29312));
    CascadeMux I__6710 (
            .O(N__29365),
            .I(N__29308));
    CascadeMux I__6709 (
            .O(N__29364),
            .I(N__29305));
    InMux I__6708 (
            .O(N__29361),
            .I(N__29302));
    InMux I__6707 (
            .O(N__29358),
            .I(N__29298));
    InMux I__6706 (
            .O(N__29357),
            .I(N__29295));
    InMux I__6705 (
            .O(N__29356),
            .I(N__29292));
    LocalMux I__6704 (
            .O(N__29353),
            .I(N__29284));
    LocalMux I__6703 (
            .O(N__29350),
            .I(N__29284));
    LocalMux I__6702 (
            .O(N__29347),
            .I(N__29284));
    LocalMux I__6701 (
            .O(N__29344),
            .I(N__29281));
    Span4Mux_v I__6700 (
            .O(N__29339),
            .I(N__29278));
    LocalMux I__6699 (
            .O(N__29336),
            .I(N__29275));
    Span4Mux_s2_v I__6698 (
            .O(N__29333),
            .I(N__29272));
    LocalMux I__6697 (
            .O(N__29330),
            .I(N__29269));
    CascadeMux I__6696 (
            .O(N__29329),
            .I(N__29266));
    InMux I__6695 (
            .O(N__29326),
            .I(N__29262));
    InMux I__6694 (
            .O(N__29323),
            .I(N__29259));
    InMux I__6693 (
            .O(N__29320),
            .I(N__29256));
    InMux I__6692 (
            .O(N__29317),
            .I(N__29253));
    InMux I__6691 (
            .O(N__29316),
            .I(N__29250));
    InMux I__6690 (
            .O(N__29315),
            .I(N__29247));
    InMux I__6689 (
            .O(N__29312),
            .I(N__29244));
    InMux I__6688 (
            .O(N__29311),
            .I(N__29241));
    InMux I__6687 (
            .O(N__29308),
            .I(N__29238));
    InMux I__6686 (
            .O(N__29305),
            .I(N__29235));
    LocalMux I__6685 (
            .O(N__29302),
            .I(N__29232));
    CascadeMux I__6684 (
            .O(N__29301),
            .I(N__29229));
    LocalMux I__6683 (
            .O(N__29298),
            .I(N__29226));
    LocalMux I__6682 (
            .O(N__29295),
            .I(N__29223));
    LocalMux I__6681 (
            .O(N__29292),
            .I(N__29220));
    InMux I__6680 (
            .O(N__29291),
            .I(N__29217));
    Span4Mux_v I__6679 (
            .O(N__29284),
            .I(N__29214));
    Span4Mux_v I__6678 (
            .O(N__29281),
            .I(N__29209));
    Span4Mux_h I__6677 (
            .O(N__29278),
            .I(N__29209));
    Span4Mux_h I__6676 (
            .O(N__29275),
            .I(N__29202));
    Span4Mux_h I__6675 (
            .O(N__29272),
            .I(N__29202));
    Span4Mux_s3_h I__6674 (
            .O(N__29269),
            .I(N__29202));
    InMux I__6673 (
            .O(N__29266),
            .I(N__29198));
    InMux I__6672 (
            .O(N__29265),
            .I(N__29195));
    LocalMux I__6671 (
            .O(N__29262),
            .I(N__29188));
    LocalMux I__6670 (
            .O(N__29259),
            .I(N__29188));
    LocalMux I__6669 (
            .O(N__29256),
            .I(N__29188));
    LocalMux I__6668 (
            .O(N__29253),
            .I(N__29185));
    LocalMux I__6667 (
            .O(N__29250),
            .I(N__29176));
    LocalMux I__6666 (
            .O(N__29247),
            .I(N__29176));
    LocalMux I__6665 (
            .O(N__29244),
            .I(N__29176));
    LocalMux I__6664 (
            .O(N__29241),
            .I(N__29176));
    LocalMux I__6663 (
            .O(N__29238),
            .I(N__29173));
    LocalMux I__6662 (
            .O(N__29235),
            .I(N__29168));
    Span4Mux_h I__6661 (
            .O(N__29232),
            .I(N__29168));
    InMux I__6660 (
            .O(N__29229),
            .I(N__29165));
    Span4Mux_s3_h I__6659 (
            .O(N__29226),
            .I(N__29158));
    Span4Mux_v I__6658 (
            .O(N__29223),
            .I(N__29158));
    Span4Mux_v I__6657 (
            .O(N__29220),
            .I(N__29158));
    LocalMux I__6656 (
            .O(N__29217),
            .I(N__29155));
    Span4Mux_h I__6655 (
            .O(N__29214),
            .I(N__29148));
    Span4Mux_h I__6654 (
            .O(N__29209),
            .I(N__29148));
    Span4Mux_v I__6653 (
            .O(N__29202),
            .I(N__29148));
    InMux I__6652 (
            .O(N__29201),
            .I(N__29145));
    LocalMux I__6651 (
            .O(N__29198),
            .I(N__29142));
    LocalMux I__6650 (
            .O(N__29195),
            .I(N__29137));
    Span12Mux_s5_h I__6649 (
            .O(N__29188),
            .I(N__29137));
    Span4Mux_s3_v I__6648 (
            .O(N__29185),
            .I(N__29132));
    Span4Mux_v I__6647 (
            .O(N__29176),
            .I(N__29132));
    Span4Mux_s3_h I__6646 (
            .O(N__29173),
            .I(N__29127));
    Span4Mux_h I__6645 (
            .O(N__29168),
            .I(N__29127));
    LocalMux I__6644 (
            .O(N__29165),
            .I(N__29122));
    Span4Mux_h I__6643 (
            .O(N__29158),
            .I(N__29122));
    Span4Mux_h I__6642 (
            .O(N__29155),
            .I(N__29117));
    Span4Mux_v I__6641 (
            .O(N__29148),
            .I(N__29117));
    LocalMux I__6640 (
            .O(N__29145),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ));
    Odrv4 I__6639 (
            .O(N__29142),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ));
    Odrv12 I__6638 (
            .O(N__29137),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ));
    Odrv4 I__6637 (
            .O(N__29132),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ));
    Odrv4 I__6636 (
            .O(N__29127),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ));
    Odrv4 I__6635 (
            .O(N__29122),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ));
    Odrv4 I__6634 (
            .O(N__29117),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ));
    CascadeMux I__6633 (
            .O(N__29102),
            .I(N__29099));
    InMux I__6632 (
            .O(N__29099),
            .I(N__29096));
    LocalMux I__6631 (
            .O(N__29096),
            .I(N__29092));
    InMux I__6630 (
            .O(N__29095),
            .I(N__29089));
    Span4Mux_s3_v I__6629 (
            .O(N__29092),
            .I(N__29084));
    LocalMux I__6628 (
            .O(N__29089),
            .I(N__29084));
    Span4Mux_v I__6627 (
            .O(N__29084),
            .I(N__29081));
    Span4Mux_h I__6626 (
            .O(N__29081),
            .I(N__29078));
    Odrv4 I__6625 (
            .O(N__29078),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_6 ));
    InMux I__6624 (
            .O(N__29075),
            .I(N__29072));
    LocalMux I__6623 (
            .O(N__29072),
            .I(N__29068));
    InMux I__6622 (
            .O(N__29071),
            .I(N__29065));
    Span4Mux_v I__6621 (
            .O(N__29068),
            .I(N__29060));
    LocalMux I__6620 (
            .O(N__29065),
            .I(N__29060));
    Span4Mux_h I__6619 (
            .O(N__29060),
            .I(N__29057));
    Odrv4 I__6618 (
            .O(N__29057),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_5 ));
    InMux I__6617 (
            .O(N__29054),
            .I(N__29048));
    InMux I__6616 (
            .O(N__29053),
            .I(N__29048));
    LocalMux I__6615 (
            .O(N__29048),
            .I(N__29045));
    Span4Mux_s3_h I__6614 (
            .O(N__29045),
            .I(N__29042));
    Span4Mux_v I__6613 (
            .O(N__29042),
            .I(N__29039));
    Odrv4 I__6612 (
            .O(N__29039),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_6 ));
    CEMux I__6611 (
            .O(N__29036),
            .I(N__29033));
    LocalMux I__6610 (
            .O(N__29033),
            .I(N__29030));
    Span4Mux_v I__6609 (
            .O(N__29030),
            .I(N__29027));
    Span4Mux_h I__6608 (
            .O(N__29027),
            .I(N__29024));
    Span4Mux_h I__6607 (
            .O(N__29024),
            .I(N__29021));
    Odrv4 I__6606 (
            .O(N__29021),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe26 ));
    CascadeMux I__6605 (
            .O(N__29018),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_7_cascade_ ));
    InMux I__6604 (
            .O(N__29015),
            .I(N__29009));
    InMux I__6603 (
            .O(N__29014),
            .I(N__29006));
    InMux I__6602 (
            .O(N__29013),
            .I(N__28994));
    InMux I__6601 (
            .O(N__29012),
            .I(N__28991));
    LocalMux I__6600 (
            .O(N__29009),
            .I(N__28988));
    LocalMux I__6599 (
            .O(N__29006),
            .I(N__28985));
    InMux I__6598 (
            .O(N__29005),
            .I(N__28982));
    InMux I__6597 (
            .O(N__29004),
            .I(N__28979));
    InMux I__6596 (
            .O(N__29003),
            .I(N__28975));
    InMux I__6595 (
            .O(N__29002),
            .I(N__28970));
    InMux I__6594 (
            .O(N__29001),
            .I(N__28965));
    InMux I__6593 (
            .O(N__29000),
            .I(N__28960));
    InMux I__6592 (
            .O(N__28999),
            .I(N__28960));
    CascadeMux I__6591 (
            .O(N__28998),
            .I(N__28951));
    InMux I__6590 (
            .O(N__28997),
            .I(N__28946));
    LocalMux I__6589 (
            .O(N__28994),
            .I(N__28921));
    LocalMux I__6588 (
            .O(N__28991),
            .I(N__28918));
    Span4Mux_s1_h I__6587 (
            .O(N__28988),
            .I(N__28909));
    Span4Mux_v I__6586 (
            .O(N__28985),
            .I(N__28909));
    LocalMux I__6585 (
            .O(N__28982),
            .I(N__28909));
    LocalMux I__6584 (
            .O(N__28979),
            .I(N__28909));
    InMux I__6583 (
            .O(N__28978),
            .I(N__28906));
    LocalMux I__6582 (
            .O(N__28975),
            .I(N__28903));
    CascadeMux I__6581 (
            .O(N__28974),
            .I(N__28900));
    InMux I__6580 (
            .O(N__28973),
            .I(N__28897));
    LocalMux I__6579 (
            .O(N__28970),
            .I(N__28894));
    InMux I__6578 (
            .O(N__28969),
            .I(N__28890));
    InMux I__6577 (
            .O(N__28968),
            .I(N__28886));
    LocalMux I__6576 (
            .O(N__28965),
            .I(N__28882));
    LocalMux I__6575 (
            .O(N__28960),
            .I(N__28879));
    InMux I__6574 (
            .O(N__28959),
            .I(N__28870));
    InMux I__6573 (
            .O(N__28958),
            .I(N__28870));
    InMux I__6572 (
            .O(N__28957),
            .I(N__28870));
    InMux I__6571 (
            .O(N__28956),
            .I(N__28870));
    InMux I__6570 (
            .O(N__28955),
            .I(N__28867));
    InMux I__6569 (
            .O(N__28954),
            .I(N__28858));
    InMux I__6568 (
            .O(N__28951),
            .I(N__28858));
    InMux I__6567 (
            .O(N__28950),
            .I(N__28858));
    InMux I__6566 (
            .O(N__28949),
            .I(N__28858));
    LocalMux I__6565 (
            .O(N__28946),
            .I(N__28855));
    InMux I__6564 (
            .O(N__28945),
            .I(N__28850));
    InMux I__6563 (
            .O(N__28944),
            .I(N__28850));
    InMux I__6562 (
            .O(N__28943),
            .I(N__28841));
    InMux I__6561 (
            .O(N__28942),
            .I(N__28841));
    InMux I__6560 (
            .O(N__28941),
            .I(N__28841));
    InMux I__6559 (
            .O(N__28940),
            .I(N__28841));
    InMux I__6558 (
            .O(N__28939),
            .I(N__28828));
    InMux I__6557 (
            .O(N__28938),
            .I(N__28828));
    InMux I__6556 (
            .O(N__28937),
            .I(N__28828));
    InMux I__6555 (
            .O(N__28936),
            .I(N__28828));
    InMux I__6554 (
            .O(N__28935),
            .I(N__28828));
    InMux I__6553 (
            .O(N__28934),
            .I(N__28828));
    InMux I__6552 (
            .O(N__28933),
            .I(N__28819));
    InMux I__6551 (
            .O(N__28932),
            .I(N__28819));
    InMux I__6550 (
            .O(N__28931),
            .I(N__28819));
    InMux I__6549 (
            .O(N__28930),
            .I(N__28819));
    InMux I__6548 (
            .O(N__28929),
            .I(N__28814));
    InMux I__6547 (
            .O(N__28928),
            .I(N__28814));
    InMux I__6546 (
            .O(N__28927),
            .I(N__28809));
    InMux I__6545 (
            .O(N__28926),
            .I(N__28809));
    InMux I__6544 (
            .O(N__28925),
            .I(N__28806));
    InMux I__6543 (
            .O(N__28924),
            .I(N__28803));
    Span4Mux_s1_h I__6542 (
            .O(N__28921),
            .I(N__28794));
    Span4Mux_v I__6541 (
            .O(N__28918),
            .I(N__28794));
    Span4Mux_v I__6540 (
            .O(N__28909),
            .I(N__28794));
    LocalMux I__6539 (
            .O(N__28906),
            .I(N__28794));
    Span4Mux_s2_h I__6538 (
            .O(N__28903),
            .I(N__28791));
    InMux I__6537 (
            .O(N__28900),
            .I(N__28788));
    LocalMux I__6536 (
            .O(N__28897),
            .I(N__28785));
    Span4Mux_v I__6535 (
            .O(N__28894),
            .I(N__28782));
    InMux I__6534 (
            .O(N__28893),
            .I(N__28775));
    LocalMux I__6533 (
            .O(N__28890),
            .I(N__28771));
    InMux I__6532 (
            .O(N__28889),
            .I(N__28768));
    LocalMux I__6531 (
            .O(N__28886),
            .I(N__28763));
    InMux I__6530 (
            .O(N__28885),
            .I(N__28760));
    Span4Mux_v I__6529 (
            .O(N__28882),
            .I(N__28749));
    Span4Mux_h I__6528 (
            .O(N__28879),
            .I(N__28749));
    LocalMux I__6527 (
            .O(N__28870),
            .I(N__28749));
    LocalMux I__6526 (
            .O(N__28867),
            .I(N__28749));
    LocalMux I__6525 (
            .O(N__28858),
            .I(N__28749));
    Span4Mux_h I__6524 (
            .O(N__28855),
            .I(N__28740));
    LocalMux I__6523 (
            .O(N__28850),
            .I(N__28740));
    LocalMux I__6522 (
            .O(N__28841),
            .I(N__28740));
    LocalMux I__6521 (
            .O(N__28828),
            .I(N__28740));
    LocalMux I__6520 (
            .O(N__28819),
            .I(N__28733));
    LocalMux I__6519 (
            .O(N__28814),
            .I(N__28733));
    LocalMux I__6518 (
            .O(N__28809),
            .I(N__28733));
    LocalMux I__6517 (
            .O(N__28806),
            .I(N__28726));
    LocalMux I__6516 (
            .O(N__28803),
            .I(N__28726));
    Span4Mux_h I__6515 (
            .O(N__28794),
            .I(N__28726));
    Sp12to4 I__6514 (
            .O(N__28791),
            .I(N__28723));
    LocalMux I__6513 (
            .O(N__28788),
            .I(N__28716));
    Span4Mux_v I__6512 (
            .O(N__28785),
            .I(N__28716));
    Span4Mux_h I__6511 (
            .O(N__28782),
            .I(N__28716));
    InMux I__6510 (
            .O(N__28781),
            .I(N__28707));
    InMux I__6509 (
            .O(N__28780),
            .I(N__28707));
    InMux I__6508 (
            .O(N__28779),
            .I(N__28707));
    InMux I__6507 (
            .O(N__28778),
            .I(N__28707));
    LocalMux I__6506 (
            .O(N__28775),
            .I(N__28704));
    InMux I__6505 (
            .O(N__28774),
            .I(N__28701));
    Span4Mux_v I__6504 (
            .O(N__28771),
            .I(N__28696));
    LocalMux I__6503 (
            .O(N__28768),
            .I(N__28696));
    InMux I__6502 (
            .O(N__28767),
            .I(N__28691));
    InMux I__6501 (
            .O(N__28766),
            .I(N__28691));
    Span4Mux_v I__6500 (
            .O(N__28763),
            .I(N__28684));
    LocalMux I__6499 (
            .O(N__28760),
            .I(N__28684));
    Span4Mux_v I__6498 (
            .O(N__28749),
            .I(N__28684));
    Span4Mux_v I__6497 (
            .O(N__28740),
            .I(N__28677));
    Span4Mux_h I__6496 (
            .O(N__28733),
            .I(N__28677));
    Span4Mux_h I__6495 (
            .O(N__28726),
            .I(N__28677));
    Odrv12 I__6494 (
            .O(N__28723),
            .I(instruction_5));
    Odrv4 I__6493 (
            .O(N__28716),
            .I(instruction_5));
    LocalMux I__6492 (
            .O(N__28707),
            .I(instruction_5));
    Odrv4 I__6491 (
            .O(N__28704),
            .I(instruction_5));
    LocalMux I__6490 (
            .O(N__28701),
            .I(instruction_5));
    Odrv4 I__6489 (
            .O(N__28696),
            .I(instruction_5));
    LocalMux I__6488 (
            .O(N__28691),
            .I(instruction_5));
    Odrv4 I__6487 (
            .O(N__28684),
            .I(instruction_5));
    Odrv4 I__6486 (
            .O(N__28677),
            .I(instruction_5));
    InMux I__6485 (
            .O(N__28658),
            .I(N__28642));
    CascadeMux I__6484 (
            .O(N__28657),
            .I(N__28634));
    InMux I__6483 (
            .O(N__28656),
            .I(N__28628));
    InMux I__6482 (
            .O(N__28655),
            .I(N__28628));
    InMux I__6481 (
            .O(N__28654),
            .I(N__28623));
    InMux I__6480 (
            .O(N__28653),
            .I(N__28623));
    InMux I__6479 (
            .O(N__28652),
            .I(N__28608));
    InMux I__6478 (
            .O(N__28651),
            .I(N__28608));
    InMux I__6477 (
            .O(N__28650),
            .I(N__28603));
    InMux I__6476 (
            .O(N__28649),
            .I(N__28603));
    InMux I__6475 (
            .O(N__28648),
            .I(N__28593));
    InMux I__6474 (
            .O(N__28647),
            .I(N__28593));
    InMux I__6473 (
            .O(N__28646),
            .I(N__28588));
    InMux I__6472 (
            .O(N__28645),
            .I(N__28588));
    LocalMux I__6471 (
            .O(N__28642),
            .I(N__28582));
    InMux I__6470 (
            .O(N__28641),
            .I(N__28577));
    InMux I__6469 (
            .O(N__28640),
            .I(N__28577));
    InMux I__6468 (
            .O(N__28639),
            .I(N__28572));
    InMux I__6467 (
            .O(N__28638),
            .I(N__28563));
    InMux I__6466 (
            .O(N__28637),
            .I(N__28563));
    InMux I__6465 (
            .O(N__28634),
            .I(N__28563));
    InMux I__6464 (
            .O(N__28633),
            .I(N__28563));
    LocalMux I__6463 (
            .O(N__28628),
            .I(N__28551));
    LocalMux I__6462 (
            .O(N__28623),
            .I(N__28551));
    InMux I__6461 (
            .O(N__28622),
            .I(N__28546));
    InMux I__6460 (
            .O(N__28621),
            .I(N__28546));
    InMux I__6459 (
            .O(N__28620),
            .I(N__28539));
    InMux I__6458 (
            .O(N__28619),
            .I(N__28539));
    InMux I__6457 (
            .O(N__28618),
            .I(N__28534));
    InMux I__6456 (
            .O(N__28617),
            .I(N__28534));
    InMux I__6455 (
            .O(N__28616),
            .I(N__28529));
    InMux I__6454 (
            .O(N__28615),
            .I(N__28529));
    InMux I__6453 (
            .O(N__28614),
            .I(N__28522));
    InMux I__6452 (
            .O(N__28613),
            .I(N__28522));
    LocalMux I__6451 (
            .O(N__28608),
            .I(N__28519));
    LocalMux I__6450 (
            .O(N__28603),
            .I(N__28516));
    InMux I__6449 (
            .O(N__28602),
            .I(N__28511));
    InMux I__6448 (
            .O(N__28601),
            .I(N__28511));
    InMux I__6447 (
            .O(N__28600),
            .I(N__28506));
    InMux I__6446 (
            .O(N__28599),
            .I(N__28506));
    InMux I__6445 (
            .O(N__28598),
            .I(N__28503));
    LocalMux I__6444 (
            .O(N__28593),
            .I(N__28498));
    LocalMux I__6443 (
            .O(N__28588),
            .I(N__28498));
    InMux I__6442 (
            .O(N__28587),
            .I(N__28495));
    InMux I__6441 (
            .O(N__28586),
            .I(N__28490));
    InMux I__6440 (
            .O(N__28585),
            .I(N__28490));
    Span4Mux_h I__6439 (
            .O(N__28582),
            .I(N__28485));
    LocalMux I__6438 (
            .O(N__28577),
            .I(N__28485));
    InMux I__6437 (
            .O(N__28576),
            .I(N__28480));
    InMux I__6436 (
            .O(N__28575),
            .I(N__28480));
    LocalMux I__6435 (
            .O(N__28572),
            .I(N__28475));
    LocalMux I__6434 (
            .O(N__28563),
            .I(N__28475));
    InMux I__6433 (
            .O(N__28562),
            .I(N__28468));
    InMux I__6432 (
            .O(N__28561),
            .I(N__28468));
    InMux I__6431 (
            .O(N__28560),
            .I(N__28468));
    InMux I__6430 (
            .O(N__28559),
            .I(N__28461));
    InMux I__6429 (
            .O(N__28558),
            .I(N__28461));
    InMux I__6428 (
            .O(N__28557),
            .I(N__28461));
    InMux I__6427 (
            .O(N__28556),
            .I(N__28458));
    Span4Mux_v I__6426 (
            .O(N__28551),
            .I(N__28453));
    LocalMux I__6425 (
            .O(N__28546),
            .I(N__28453));
    InMux I__6424 (
            .O(N__28545),
            .I(N__28448));
    InMux I__6423 (
            .O(N__28544),
            .I(N__28448));
    LocalMux I__6422 (
            .O(N__28539),
            .I(N__28443));
    LocalMux I__6421 (
            .O(N__28534),
            .I(N__28443));
    LocalMux I__6420 (
            .O(N__28529),
            .I(N__28437));
    InMux I__6419 (
            .O(N__28528),
            .I(N__28432));
    InMux I__6418 (
            .O(N__28527),
            .I(N__28432));
    LocalMux I__6417 (
            .O(N__28522),
            .I(N__28429));
    Span4Mux_v I__6416 (
            .O(N__28519),
            .I(N__28420));
    Span4Mux_v I__6415 (
            .O(N__28516),
            .I(N__28420));
    LocalMux I__6414 (
            .O(N__28511),
            .I(N__28415));
    LocalMux I__6413 (
            .O(N__28506),
            .I(N__28415));
    LocalMux I__6412 (
            .O(N__28503),
            .I(N__28406));
    Span4Mux_v I__6411 (
            .O(N__28498),
            .I(N__28406));
    LocalMux I__6410 (
            .O(N__28495),
            .I(N__28406));
    LocalMux I__6409 (
            .O(N__28490),
            .I(N__28406));
    Span4Mux_s3_h I__6408 (
            .O(N__28485),
            .I(N__28401));
    LocalMux I__6407 (
            .O(N__28480),
            .I(N__28401));
    Span4Mux_v I__6406 (
            .O(N__28475),
            .I(N__28392));
    LocalMux I__6405 (
            .O(N__28468),
            .I(N__28392));
    LocalMux I__6404 (
            .O(N__28461),
            .I(N__28392));
    LocalMux I__6403 (
            .O(N__28458),
            .I(N__28392));
    Span4Mux_h I__6402 (
            .O(N__28453),
            .I(N__28385));
    LocalMux I__6401 (
            .O(N__28448),
            .I(N__28385));
    Span4Mux_v I__6400 (
            .O(N__28443),
            .I(N__28385));
    InMux I__6399 (
            .O(N__28442),
            .I(N__28378));
    InMux I__6398 (
            .O(N__28441),
            .I(N__28378));
    InMux I__6397 (
            .O(N__28440),
            .I(N__28378));
    Span4Mux_s1_h I__6396 (
            .O(N__28437),
            .I(N__28373));
    LocalMux I__6395 (
            .O(N__28432),
            .I(N__28373));
    Span4Mux_v I__6394 (
            .O(N__28429),
            .I(N__28370));
    InMux I__6393 (
            .O(N__28428),
            .I(N__28365));
    InMux I__6392 (
            .O(N__28427),
            .I(N__28365));
    InMux I__6391 (
            .O(N__28426),
            .I(N__28360));
    InMux I__6390 (
            .O(N__28425),
            .I(N__28360));
    Span4Mux_h I__6389 (
            .O(N__28420),
            .I(N__28353));
    Span4Mux_v I__6388 (
            .O(N__28415),
            .I(N__28353));
    Span4Mux_v I__6387 (
            .O(N__28406),
            .I(N__28353));
    Span4Mux_v I__6386 (
            .O(N__28401),
            .I(N__28346));
    Span4Mux_v I__6385 (
            .O(N__28392),
            .I(N__28346));
    Span4Mux_h I__6384 (
            .O(N__28385),
            .I(N__28346));
    LocalMux I__6383 (
            .O(N__28378),
            .I(instruction_6));
    Odrv4 I__6382 (
            .O(N__28373),
            .I(instruction_6));
    Odrv4 I__6381 (
            .O(N__28370),
            .I(instruction_6));
    LocalMux I__6380 (
            .O(N__28365),
            .I(instruction_6));
    LocalMux I__6379 (
            .O(N__28360),
            .I(instruction_6));
    Odrv4 I__6378 (
            .O(N__28353),
            .I(instruction_6));
    Odrv4 I__6377 (
            .O(N__28346),
            .I(instruction_6));
    InMux I__6376 (
            .O(N__28331),
            .I(N__28328));
    LocalMux I__6375 (
            .O(N__28328),
            .I(N__28325));
    Span4Mux_s0_h I__6374 (
            .O(N__28325),
            .I(N__28322));
    Odrv4 I__6373 (
            .O(N__28322),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_7 ));
    CascadeMux I__6372 (
            .O(N__28319),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_7_cascade_ ));
    InMux I__6371 (
            .O(N__28316),
            .I(N__28313));
    LocalMux I__6370 (
            .O(N__28313),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_7 ));
    InMux I__6369 (
            .O(N__28310),
            .I(N__28307));
    LocalMux I__6368 (
            .O(N__28307),
            .I(N__28304));
    Span4Mux_v I__6367 (
            .O(N__28304),
            .I(N__28301));
    Span4Mux_h I__6366 (
            .O(N__28301),
            .I(N__28298));
    Span4Mux_h I__6365 (
            .O(N__28298),
            .I(N__28295));
    Odrv4 I__6364 (
            .O(N__28295),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_7 ));
    InMux I__6363 (
            .O(N__28292),
            .I(N__28288));
    InMux I__6362 (
            .O(N__28291),
            .I(N__28285));
    LocalMux I__6361 (
            .O(N__28288),
            .I(N__28280));
    LocalMux I__6360 (
            .O(N__28285),
            .I(N__28280));
    Odrv4 I__6359 (
            .O(N__28280),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_7 ));
    CascadeMux I__6358 (
            .O(N__28277),
            .I(N__28274));
    InMux I__6357 (
            .O(N__28274),
            .I(N__28268));
    InMux I__6356 (
            .O(N__28273),
            .I(N__28268));
    LocalMux I__6355 (
            .O(N__28268),
            .I(N__28265));
    Odrv12 I__6354 (
            .O(N__28265),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_7 ));
    CascadeMux I__6353 (
            .O(N__28262),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_7_cascade_ ));
    InMux I__6352 (
            .O(N__28259),
            .I(N__28256));
    LocalMux I__6351 (
            .O(N__28256),
            .I(N__28253));
    Span4Mux_h I__6350 (
            .O(N__28253),
            .I(N__28250));
    Span4Mux_h I__6349 (
            .O(N__28250),
            .I(N__28247));
    Odrv4 I__6348 (
            .O(N__28247),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI0NMM1_7 ));
    CascadeMux I__6347 (
            .O(N__28244),
            .I(N__28241));
    InMux I__6346 (
            .O(N__28241),
            .I(N__28237));
    CascadeMux I__6345 (
            .O(N__28240),
            .I(N__28234));
    LocalMux I__6344 (
            .O(N__28237),
            .I(N__28231));
    InMux I__6343 (
            .O(N__28234),
            .I(N__28228));
    Span4Mux_h I__6342 (
            .O(N__28231),
            .I(N__28225));
    LocalMux I__6341 (
            .O(N__28228),
            .I(N__28222));
    Odrv4 I__6340 (
            .O(N__28225),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4 ));
    Odrv4 I__6339 (
            .O(N__28222),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4 ));
    CascadeMux I__6338 (
            .O(N__28217),
            .I(N__28213));
    InMux I__6337 (
            .O(N__28216),
            .I(N__28208));
    InMux I__6336 (
            .O(N__28213),
            .I(N__28208));
    LocalMux I__6335 (
            .O(N__28208),
            .I(N__28205));
    Span4Mux_v I__6334 (
            .O(N__28205),
            .I(N__28202));
    Odrv4 I__6333 (
            .O(N__28202),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_5 ));
    InMux I__6332 (
            .O(N__28199),
            .I(N__28195));
    InMux I__6331 (
            .O(N__28198),
            .I(N__28192));
    LocalMux I__6330 (
            .O(N__28195),
            .I(N__28187));
    LocalMux I__6329 (
            .O(N__28192),
            .I(N__28187));
    Span4Mux_h I__6328 (
            .O(N__28187),
            .I(N__28184));
    Odrv4 I__6327 (
            .O(N__28184),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_6 ));
    CEMux I__6326 (
            .O(N__28181),
            .I(N__28178));
    LocalMux I__6325 (
            .O(N__28178),
            .I(N__28175));
    Span4Mux_s3_h I__6324 (
            .O(N__28175),
            .I(N__28172));
    Span4Mux_v I__6323 (
            .O(N__28172),
            .I(N__28169));
    Span4Mux_h I__6322 (
            .O(N__28169),
            .I(N__28166));
    Odrv4 I__6321 (
            .O(N__28166),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe25 ));
    InMux I__6320 (
            .O(N__28163),
            .I(N__28160));
    LocalMux I__6319 (
            .O(N__28160),
            .I(N__28156));
    InMux I__6318 (
            .O(N__28159),
            .I(N__28153));
    Span4Mux_h I__6317 (
            .O(N__28156),
            .I(N__28150));
    LocalMux I__6316 (
            .O(N__28153),
            .I(N__28147));
    Odrv4 I__6315 (
            .O(N__28150),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0 ));
    Odrv12 I__6314 (
            .O(N__28147),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0 ));
    InMux I__6313 (
            .O(N__28142),
            .I(N__28136));
    InMux I__6312 (
            .O(N__28141),
            .I(N__28136));
    LocalMux I__6311 (
            .O(N__28136),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_1 ));
    InMux I__6310 (
            .O(N__28133),
            .I(N__28130));
    LocalMux I__6309 (
            .O(N__28130),
            .I(N__28126));
    CascadeMux I__6308 (
            .O(N__28129),
            .I(N__28123));
    Span4Mux_v I__6307 (
            .O(N__28126),
            .I(N__28120));
    InMux I__6306 (
            .O(N__28123),
            .I(N__28117));
    Odrv4 I__6305 (
            .O(N__28120),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2 ));
    LocalMux I__6304 (
            .O(N__28117),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2 ));
    InMux I__6303 (
            .O(N__28112),
            .I(N__28109));
    LocalMux I__6302 (
            .O(N__28109),
            .I(N__28105));
    InMux I__6301 (
            .O(N__28108),
            .I(N__28102));
    Span4Mux_v I__6300 (
            .O(N__28105),
            .I(N__28099));
    LocalMux I__6299 (
            .O(N__28102),
            .I(N__28096));
    Odrv4 I__6298 (
            .O(N__28099),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3 ));
    Odrv4 I__6297 (
            .O(N__28096),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3 ));
    InMux I__6296 (
            .O(N__28091),
            .I(N__28088));
    LocalMux I__6295 (
            .O(N__28088),
            .I(N__28085));
    Span4Mux_v I__6294 (
            .O(N__28085),
            .I(N__28081));
    InMux I__6293 (
            .O(N__28084),
            .I(N__28078));
    Span4Mux_h I__6292 (
            .O(N__28081),
            .I(N__28075));
    LocalMux I__6291 (
            .O(N__28078),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4 ));
    Odrv4 I__6290 (
            .O(N__28075),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4 ));
    InMux I__6289 (
            .O(N__28070),
            .I(N__28064));
    InMux I__6288 (
            .O(N__28069),
            .I(N__28064));
    LocalMux I__6287 (
            .O(N__28064),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_3 ));
    InMux I__6286 (
            .O(N__28061),
            .I(N__28057));
    InMux I__6285 (
            .O(N__28060),
            .I(N__28054));
    LocalMux I__6284 (
            .O(N__28057),
            .I(N__28051));
    LocalMux I__6283 (
            .O(N__28054),
            .I(N__28048));
    Span4Mux_v I__6282 (
            .O(N__28051),
            .I(N__28045));
    Span4Mux_v I__6281 (
            .O(N__28048),
            .I(N__28042));
    Odrv4 I__6280 (
            .O(N__28045),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4 ));
    Odrv4 I__6279 (
            .O(N__28042),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4 ));
    InMux I__6278 (
            .O(N__28037),
            .I(N__28031));
    InMux I__6277 (
            .O(N__28036),
            .I(N__28031));
    LocalMux I__6276 (
            .O(N__28031),
            .I(N__28028));
    Span4Mux_h I__6275 (
            .O(N__28028),
            .I(N__28025));
    Odrv4 I__6274 (
            .O(N__28025),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_5 ));
    CascadeMux I__6273 (
            .O(N__28022),
            .I(N__28019));
    InMux I__6272 (
            .O(N__28019),
            .I(N__28013));
    InMux I__6271 (
            .O(N__28018),
            .I(N__28013));
    LocalMux I__6270 (
            .O(N__28013),
            .I(N__28010));
    Span4Mux_h I__6269 (
            .O(N__28010),
            .I(N__28007));
    Odrv4 I__6268 (
            .O(N__28007),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_6 ));
    CEMux I__6267 (
            .O(N__28004),
            .I(N__28001));
    LocalMux I__6266 (
            .O(N__28001),
            .I(N__27998));
    Span4Mux_s0_h I__6265 (
            .O(N__27998),
            .I(N__27995));
    Span4Mux_h I__6264 (
            .O(N__27995),
            .I(N__27992));
    Odrv4 I__6263 (
            .O(N__27992),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe24 ));
    CascadeMux I__6262 (
            .O(N__27989),
            .I(N__27985));
    InMux I__6261 (
            .O(N__27988),
            .I(N__27980));
    InMux I__6260 (
            .O(N__27985),
            .I(N__27980));
    LocalMux I__6259 (
            .O(N__27980),
            .I(N__27977));
    Span4Mux_h I__6258 (
            .O(N__27977),
            .I(N__27974));
    Odrv4 I__6257 (
            .O(N__27974),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_0 ));
    CascadeMux I__6256 (
            .O(N__27971),
            .I(N__27968));
    InMux I__6255 (
            .O(N__27968),
            .I(N__27964));
    CascadeMux I__6254 (
            .O(N__27967),
            .I(N__27961));
    LocalMux I__6253 (
            .O(N__27964),
            .I(N__27958));
    InMux I__6252 (
            .O(N__27961),
            .I(N__27955));
    Odrv4 I__6251 (
            .O(N__27958),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1 ));
    LocalMux I__6250 (
            .O(N__27955),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1 ));
    InMux I__6249 (
            .O(N__27950),
            .I(N__27944));
    InMux I__6248 (
            .O(N__27949),
            .I(N__27944));
    LocalMux I__6247 (
            .O(N__27944),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_2 ));
    InMux I__6246 (
            .O(N__27941),
            .I(N__27935));
    InMux I__6245 (
            .O(N__27940),
            .I(N__27935));
    LocalMux I__6244 (
            .O(N__27935),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_3 ));
    InMux I__6243 (
            .O(N__27932),
            .I(N__27929));
    LocalMux I__6242 (
            .O(N__27929),
            .I(N__27925));
    InMux I__6241 (
            .O(N__27928),
            .I(N__27922));
    Span4Mux_v I__6240 (
            .O(N__27925),
            .I(N__27917));
    LocalMux I__6239 (
            .O(N__27922),
            .I(N__27917));
    Span4Mux_v I__6238 (
            .O(N__27917),
            .I(N__27914));
    Odrv4 I__6237 (
            .O(N__27914),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_3 ));
    CascadeMux I__6236 (
            .O(N__27911),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_3_cascade_ ));
    InMux I__6235 (
            .O(N__27908),
            .I(N__27904));
    InMux I__6234 (
            .O(N__27907),
            .I(N__27901));
    LocalMux I__6233 (
            .O(N__27904),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3 ));
    LocalMux I__6232 (
            .O(N__27901),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3 ));
    InMux I__6231 (
            .O(N__27896),
            .I(N__27893));
    LocalMux I__6230 (
            .O(N__27893),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIKIUU1_3 ));
    CascadeMux I__6229 (
            .O(N__27890),
            .I(N__27887));
    InMux I__6228 (
            .O(N__27887),
            .I(N__27883));
    InMux I__6227 (
            .O(N__27886),
            .I(N__27880));
    LocalMux I__6226 (
            .O(N__27883),
            .I(N__27877));
    LocalMux I__6225 (
            .O(N__27880),
            .I(N__27874));
    Span4Mux_v I__6224 (
            .O(N__27877),
            .I(N__27869));
    Span4Mux_v I__6223 (
            .O(N__27874),
            .I(N__27869));
    Odrv4 I__6222 (
            .O(N__27869),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_3 ));
    InMux I__6221 (
            .O(N__27866),
            .I(N__27862));
    InMux I__6220 (
            .O(N__27865),
            .I(N__27859));
    LocalMux I__6219 (
            .O(N__27862),
            .I(N__27856));
    LocalMux I__6218 (
            .O(N__27859),
            .I(N__27853));
    Span4Mux_s3_h I__6217 (
            .O(N__27856),
            .I(N__27850));
    Span4Mux_s2_h I__6216 (
            .O(N__27853),
            .I(N__27847));
    Odrv4 I__6215 (
            .O(N__27850),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3 ));
    Odrv4 I__6214 (
            .O(N__27847),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3 ));
    InMux I__6213 (
            .O(N__27842),
            .I(N__27839));
    LocalMux I__6212 (
            .O(N__27839),
            .I(N__27836));
    Odrv4 I__6211 (
            .O(N__27836),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_3 ));
    CascadeMux I__6210 (
            .O(N__27833),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_3_cascade_ ));
    CascadeMux I__6209 (
            .O(N__27830),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_3_cascade_ ));
    InMux I__6208 (
            .O(N__27827),
            .I(N__27824));
    LocalMux I__6207 (
            .O(N__27824),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_3 ));
    InMux I__6206 (
            .O(N__27821),
            .I(N__27818));
    LocalMux I__6205 (
            .O(N__27818),
            .I(N__27815));
    Span4Mux_h I__6204 (
            .O(N__27815),
            .I(N__27812));
    Odrv4 I__6203 (
            .O(N__27812),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_3 ));
    InMux I__6202 (
            .O(N__27809),
            .I(N__27805));
    InMux I__6201 (
            .O(N__27808),
            .I(N__27802));
    LocalMux I__6200 (
            .O(N__27805),
            .I(N__27799));
    LocalMux I__6199 (
            .O(N__27802),
            .I(N__27796));
    Span12Mux_s1_h I__6198 (
            .O(N__27799),
            .I(N__27791));
    Span12Mux_s7_v I__6197 (
            .O(N__27796),
            .I(N__27791));
    Odrv12 I__6196 (
            .O(N__27791),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_2 ));
    CEMux I__6195 (
            .O(N__27788),
            .I(N__27785));
    LocalMux I__6194 (
            .O(N__27785),
            .I(N__27782));
    Span4Mux_v I__6193 (
            .O(N__27782),
            .I(N__27778));
    CEMux I__6192 (
            .O(N__27781),
            .I(N__27775));
    Span4Mux_h I__6191 (
            .O(N__27778),
            .I(N__27771));
    LocalMux I__6190 (
            .O(N__27775),
            .I(N__27768));
    CEMux I__6189 (
            .O(N__27774),
            .I(N__27765));
    Span4Mux_v I__6188 (
            .O(N__27771),
            .I(N__27762));
    Span4Mux_h I__6187 (
            .O(N__27768),
            .I(N__27759));
    LocalMux I__6186 (
            .O(N__27765),
            .I(N__27756));
    Odrv4 I__6185 (
            .O(N__27762),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31 ));
    Odrv4 I__6184 (
            .O(N__27759),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31 ));
    Odrv12 I__6183 (
            .O(N__27756),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31 ));
    InMux I__6182 (
            .O(N__27749),
            .I(N__27743));
    InMux I__6181 (
            .O(N__27748),
            .I(N__27743));
    LocalMux I__6180 (
            .O(N__27743),
            .I(N__27740));
    Span4Mux_h I__6179 (
            .O(N__27740),
            .I(N__27737));
    Odrv4 I__6178 (
            .O(N__27737),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_0 ));
    InMux I__6177 (
            .O(N__27734),
            .I(N__27731));
    LocalMux I__6176 (
            .O(N__27731),
            .I(N__27728));
    Span4Mux_v I__6175 (
            .O(N__27728),
            .I(N__27724));
    InMux I__6174 (
            .O(N__27727),
            .I(N__27721));
    Odrv4 I__6173 (
            .O(N__27724),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1 ));
    LocalMux I__6172 (
            .O(N__27721),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1 ));
    InMux I__6171 (
            .O(N__27716),
            .I(N__27710));
    InMux I__6170 (
            .O(N__27715),
            .I(N__27710));
    LocalMux I__6169 (
            .O(N__27710),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_2 ));
    InMux I__6168 (
            .O(N__27707),
            .I(N__27703));
    InMux I__6167 (
            .O(N__27706),
            .I(N__27700));
    LocalMux I__6166 (
            .O(N__27703),
            .I(N__27697));
    LocalMux I__6165 (
            .O(N__27700),
            .I(N__27692));
    Span4Mux_h I__6164 (
            .O(N__27697),
            .I(N__27692));
    Span4Mux_h I__6163 (
            .O(N__27692),
            .I(N__27689));
    Odrv4 I__6162 (
            .O(N__27689),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_4 ));
    CEMux I__6161 (
            .O(N__27686),
            .I(N__27683));
    LocalMux I__6160 (
            .O(N__27683),
            .I(N__27680));
    Span4Mux_v I__6159 (
            .O(N__27680),
            .I(N__27676));
    CEMux I__6158 (
            .O(N__27679),
            .I(N__27673));
    Span4Mux_s0_h I__6157 (
            .O(N__27676),
            .I(N__27670));
    LocalMux I__6156 (
            .O(N__27673),
            .I(N__27667));
    Span4Mux_h I__6155 (
            .O(N__27670),
            .I(N__27664));
    Span4Mux_s1_v I__6154 (
            .O(N__27667),
            .I(N__27661));
    Span4Mux_h I__6153 (
            .O(N__27664),
            .I(N__27658));
    Span4Mux_h I__6152 (
            .O(N__27661),
            .I(N__27655));
    Span4Mux_s3_h I__6151 (
            .O(N__27658),
            .I(N__27652));
    Odrv4 I__6150 (
            .O(N__27655),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18 ));
    Odrv4 I__6149 (
            .O(N__27652),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18 ));
    CascadeMux I__6148 (
            .O(N__27647),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_3_cascade_ ));
    CascadeMux I__6147 (
            .O(N__27644),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI06K32_3_cascade_ ));
    InMux I__6146 (
            .O(N__27641),
            .I(N__27637));
    InMux I__6145 (
            .O(N__27640),
            .I(N__27633));
    LocalMux I__6144 (
            .O(N__27637),
            .I(N__27625));
    InMux I__6143 (
            .O(N__27636),
            .I(N__27621));
    LocalMux I__6142 (
            .O(N__27633),
            .I(N__27618));
    InMux I__6141 (
            .O(N__27632),
            .I(N__27615));
    InMux I__6140 (
            .O(N__27631),
            .I(N__27612));
    InMux I__6139 (
            .O(N__27630),
            .I(N__27606));
    InMux I__6138 (
            .O(N__27629),
            .I(N__27602));
    InMux I__6137 (
            .O(N__27628),
            .I(N__27599));
    Span4Mux_v I__6136 (
            .O(N__27625),
            .I(N__27596));
    CascadeMux I__6135 (
            .O(N__27624),
            .I(N__27591));
    LocalMux I__6134 (
            .O(N__27621),
            .I(N__27587));
    Span4Mux_v I__6133 (
            .O(N__27618),
            .I(N__27582));
    LocalMux I__6132 (
            .O(N__27615),
            .I(N__27582));
    LocalMux I__6131 (
            .O(N__27612),
            .I(N__27579));
    InMux I__6130 (
            .O(N__27611),
            .I(N__27574));
    InMux I__6129 (
            .O(N__27610),
            .I(N__27574));
    InMux I__6128 (
            .O(N__27609),
            .I(N__27571));
    LocalMux I__6127 (
            .O(N__27606),
            .I(N__27568));
    InMux I__6126 (
            .O(N__27605),
            .I(N__27565));
    LocalMux I__6125 (
            .O(N__27602),
            .I(N__27559));
    LocalMux I__6124 (
            .O(N__27599),
            .I(N__27559));
    Span4Mux_v I__6123 (
            .O(N__27596),
            .I(N__27556));
    InMux I__6122 (
            .O(N__27595),
            .I(N__27551));
    InMux I__6121 (
            .O(N__27594),
            .I(N__27551));
    InMux I__6120 (
            .O(N__27591),
            .I(N__27545));
    InMux I__6119 (
            .O(N__27590),
            .I(N__27545));
    Span4Mux_s2_h I__6118 (
            .O(N__27587),
            .I(N__27542));
    Span4Mux_h I__6117 (
            .O(N__27582),
            .I(N__27536));
    Span4Mux_h I__6116 (
            .O(N__27579),
            .I(N__27533));
    LocalMux I__6115 (
            .O(N__27574),
            .I(N__27524));
    LocalMux I__6114 (
            .O(N__27571),
            .I(N__27524));
    Span4Mux_h I__6113 (
            .O(N__27568),
            .I(N__27524));
    LocalMux I__6112 (
            .O(N__27565),
            .I(N__27524));
    InMux I__6111 (
            .O(N__27564),
            .I(N__27521));
    Span4Mux_h I__6110 (
            .O(N__27559),
            .I(N__27518));
    Span4Mux_h I__6109 (
            .O(N__27556),
            .I(N__27513));
    LocalMux I__6108 (
            .O(N__27551),
            .I(N__27513));
    InMux I__6107 (
            .O(N__27550),
            .I(N__27510));
    LocalMux I__6106 (
            .O(N__27545),
            .I(N__27505));
    Span4Mux_h I__6105 (
            .O(N__27542),
            .I(N__27505));
    InMux I__6104 (
            .O(N__27541),
            .I(N__27502));
    InMux I__6103 (
            .O(N__27540),
            .I(N__27499));
    InMux I__6102 (
            .O(N__27539),
            .I(N__27496));
    Span4Mux_v I__6101 (
            .O(N__27536),
            .I(N__27493));
    Span4Mux_v I__6100 (
            .O(N__27533),
            .I(N__27486));
    Span4Mux_v I__6099 (
            .O(N__27524),
            .I(N__27486));
    LocalMux I__6098 (
            .O(N__27521),
            .I(N__27486));
    Span4Mux_v I__6097 (
            .O(N__27518),
            .I(N__27479));
    Span4Mux_h I__6096 (
            .O(N__27513),
            .I(N__27479));
    LocalMux I__6095 (
            .O(N__27510),
            .I(N__27479));
    Span4Mux_h I__6094 (
            .O(N__27505),
            .I(N__27472));
    LocalMux I__6093 (
            .O(N__27502),
            .I(N__27472));
    LocalMux I__6092 (
            .O(N__27499),
            .I(N__27472));
    LocalMux I__6091 (
            .O(N__27496),
            .I(instruction_10));
    Odrv4 I__6090 (
            .O(N__27493),
            .I(instruction_10));
    Odrv4 I__6089 (
            .O(N__27486),
            .I(instruction_10));
    Odrv4 I__6088 (
            .O(N__27479),
            .I(instruction_10));
    Odrv4 I__6087 (
            .O(N__27472),
            .I(instruction_10));
    CascadeMux I__6086 (
            .O(N__27461),
            .I(N__27457));
    CascadeMux I__6085 (
            .O(N__27460),
            .I(N__27436));
    InMux I__6084 (
            .O(N__27457),
            .I(N__27425));
    InMux I__6083 (
            .O(N__27456),
            .I(N__27410));
    InMux I__6082 (
            .O(N__27455),
            .I(N__27410));
    InMux I__6081 (
            .O(N__27454),
            .I(N__27410));
    InMux I__6080 (
            .O(N__27453),
            .I(N__27410));
    InMux I__6079 (
            .O(N__27452),
            .I(N__27410));
    InMux I__6078 (
            .O(N__27451),
            .I(N__27410));
    InMux I__6077 (
            .O(N__27450),
            .I(N__27410));
    InMux I__6076 (
            .O(N__27449),
            .I(N__27395));
    InMux I__6075 (
            .O(N__27448),
            .I(N__27395));
    InMux I__6074 (
            .O(N__27447),
            .I(N__27395));
    InMux I__6073 (
            .O(N__27446),
            .I(N__27395));
    InMux I__6072 (
            .O(N__27445),
            .I(N__27395));
    InMux I__6071 (
            .O(N__27444),
            .I(N__27395));
    InMux I__6070 (
            .O(N__27443),
            .I(N__27395));
    InMux I__6069 (
            .O(N__27442),
            .I(N__27381));
    InMux I__6068 (
            .O(N__27441),
            .I(N__27374));
    InMux I__6067 (
            .O(N__27440),
            .I(N__27374));
    InMux I__6066 (
            .O(N__27439),
            .I(N__27374));
    InMux I__6065 (
            .O(N__27436),
            .I(N__27371));
    InMux I__6064 (
            .O(N__27435),
            .I(N__27354));
    InMux I__6063 (
            .O(N__27434),
            .I(N__27354));
    InMux I__6062 (
            .O(N__27433),
            .I(N__27354));
    InMux I__6061 (
            .O(N__27432),
            .I(N__27354));
    InMux I__6060 (
            .O(N__27431),
            .I(N__27354));
    InMux I__6059 (
            .O(N__27430),
            .I(N__27354));
    InMux I__6058 (
            .O(N__27429),
            .I(N__27354));
    InMux I__6057 (
            .O(N__27428),
            .I(N__27354));
    LocalMux I__6056 (
            .O(N__27425),
            .I(N__27347));
    LocalMux I__6055 (
            .O(N__27410),
            .I(N__27347));
    LocalMux I__6054 (
            .O(N__27395),
            .I(N__27347));
    InMux I__6053 (
            .O(N__27394),
            .I(N__27332));
    InMux I__6052 (
            .O(N__27393),
            .I(N__27332));
    InMux I__6051 (
            .O(N__27392),
            .I(N__27332));
    InMux I__6050 (
            .O(N__27391),
            .I(N__27332));
    InMux I__6049 (
            .O(N__27390),
            .I(N__27332));
    InMux I__6048 (
            .O(N__27389),
            .I(N__27332));
    InMux I__6047 (
            .O(N__27388),
            .I(N__27332));
    InMux I__6046 (
            .O(N__27387),
            .I(N__27327));
    InMux I__6045 (
            .O(N__27386),
            .I(N__27327));
    InMux I__6044 (
            .O(N__27385),
            .I(N__27322));
    InMux I__6043 (
            .O(N__27384),
            .I(N__27322));
    LocalMux I__6042 (
            .O(N__27381),
            .I(N__27317));
    LocalMux I__6041 (
            .O(N__27374),
            .I(N__27309));
    LocalMux I__6040 (
            .O(N__27371),
            .I(N__27298));
    LocalMux I__6039 (
            .O(N__27354),
            .I(N__27298));
    Span4Mux_v I__6038 (
            .O(N__27347),
            .I(N__27298));
    LocalMux I__6037 (
            .O(N__27332),
            .I(N__27298));
    LocalMux I__6036 (
            .O(N__27327),
            .I(N__27298));
    LocalMux I__6035 (
            .O(N__27322),
            .I(N__27295));
    InMux I__6034 (
            .O(N__27321),
            .I(N__27290));
    InMux I__6033 (
            .O(N__27320),
            .I(N__27290));
    Span4Mux_v I__6032 (
            .O(N__27317),
            .I(N__27282));
    InMux I__6031 (
            .O(N__27316),
            .I(N__27279));
    InMux I__6030 (
            .O(N__27315),
            .I(N__27268));
    InMux I__6029 (
            .O(N__27314),
            .I(N__27268));
    InMux I__6028 (
            .O(N__27313),
            .I(N__27263));
    InMux I__6027 (
            .O(N__27312),
            .I(N__27263));
    Span4Mux_h I__6026 (
            .O(N__27309),
            .I(N__27260));
    Span4Mux_h I__6025 (
            .O(N__27298),
            .I(N__27253));
    Span4Mux_s3_v I__6024 (
            .O(N__27295),
            .I(N__27253));
    LocalMux I__6023 (
            .O(N__27290),
            .I(N__27253));
    InMux I__6022 (
            .O(N__27289),
            .I(N__27248));
    InMux I__6021 (
            .O(N__27288),
            .I(N__27245));
    InMux I__6020 (
            .O(N__27287),
            .I(N__27242));
    InMux I__6019 (
            .O(N__27286),
            .I(N__27239));
    InMux I__6018 (
            .O(N__27285),
            .I(N__27236));
    Span4Mux_s1_h I__6017 (
            .O(N__27282),
            .I(N__27231));
    LocalMux I__6016 (
            .O(N__27279),
            .I(N__27231));
    InMux I__6015 (
            .O(N__27278),
            .I(N__27226));
    InMux I__6014 (
            .O(N__27277),
            .I(N__27226));
    InMux I__6013 (
            .O(N__27276),
            .I(N__27217));
    InMux I__6012 (
            .O(N__27275),
            .I(N__27217));
    InMux I__6011 (
            .O(N__27274),
            .I(N__27217));
    InMux I__6010 (
            .O(N__27273),
            .I(N__27217));
    LocalMux I__6009 (
            .O(N__27268),
            .I(N__27212));
    LocalMux I__6008 (
            .O(N__27263),
            .I(N__27212));
    Span4Mux_h I__6007 (
            .O(N__27260),
            .I(N__27207));
    Span4Mux_v I__6006 (
            .O(N__27253),
            .I(N__27207));
    InMux I__6005 (
            .O(N__27252),
            .I(N__27200));
    InMux I__6004 (
            .O(N__27251),
            .I(N__27200));
    LocalMux I__6003 (
            .O(N__27248),
            .I(N__27193));
    LocalMux I__6002 (
            .O(N__27245),
            .I(N__27193));
    LocalMux I__6001 (
            .O(N__27242),
            .I(N__27193));
    LocalMux I__6000 (
            .O(N__27239),
            .I(N__27188));
    LocalMux I__5999 (
            .O(N__27236),
            .I(N__27183));
    Span4Mux_h I__5998 (
            .O(N__27231),
            .I(N__27178));
    LocalMux I__5997 (
            .O(N__27226),
            .I(N__27178));
    LocalMux I__5996 (
            .O(N__27217),
            .I(N__27173));
    Span4Mux_v I__5995 (
            .O(N__27212),
            .I(N__27173));
    IoSpan4Mux I__5994 (
            .O(N__27207),
            .I(N__27170));
    InMux I__5993 (
            .O(N__27206),
            .I(N__27165));
    InMux I__5992 (
            .O(N__27205),
            .I(N__27165));
    LocalMux I__5991 (
            .O(N__27200),
            .I(N__27160));
    Span4Mux_v I__5990 (
            .O(N__27193),
            .I(N__27160));
    InMux I__5989 (
            .O(N__27192),
            .I(N__27155));
    InMux I__5988 (
            .O(N__27191),
            .I(N__27155));
    Span12Mux_s9_h I__5987 (
            .O(N__27188),
            .I(N__27152));
    InMux I__5986 (
            .O(N__27187),
            .I(N__27147));
    InMux I__5985 (
            .O(N__27186),
            .I(N__27147));
    Span4Mux_h I__5984 (
            .O(N__27183),
            .I(N__27142));
    Span4Mux_h I__5983 (
            .O(N__27178),
            .I(N__27142));
    Span4Mux_h I__5982 (
            .O(N__27173),
            .I(N__27131));
    Span4Mux_s1_h I__5981 (
            .O(N__27170),
            .I(N__27131));
    LocalMux I__5980 (
            .O(N__27165),
            .I(N__27131));
    Span4Mux_h I__5979 (
            .O(N__27160),
            .I(N__27131));
    LocalMux I__5978 (
            .O(N__27155),
            .I(N__27131));
    Odrv12 I__5977 (
            .O(N__27152),
            .I(instruction_11));
    LocalMux I__5976 (
            .O(N__27147),
            .I(instruction_11));
    Odrv4 I__5975 (
            .O(N__27142),
            .I(instruction_11));
    Odrv4 I__5974 (
            .O(N__27131),
            .I(instruction_11));
    InMux I__5973 (
            .O(N__27122),
            .I(N__27119));
    LocalMux I__5972 (
            .O(N__27119),
            .I(N__27116));
    Odrv12 I__5971 (
            .O(N__27116),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIE0IQ1_3 ));
    CascadeMux I__5970 (
            .O(N__27113),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_3_cascade_ ));
    InMux I__5969 (
            .O(N__27110),
            .I(N__27107));
    LocalMux I__5968 (
            .O(N__27107),
            .I(N__27104));
    Span4Mux_v I__5967 (
            .O(N__27104),
            .I(N__27101));
    Span4Mux_h I__5966 (
            .O(N__27101),
            .I(N__27098));
    Odrv4 I__5965 (
            .O(N__27098),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV1BI8_3 ));
    InMux I__5964 (
            .O(N__27095),
            .I(N__27091));
    InMux I__5963 (
            .O(N__27094),
            .I(N__27088));
    LocalMux I__5962 (
            .O(N__27091),
            .I(N__27085));
    LocalMux I__5961 (
            .O(N__27088),
            .I(N__27082));
    Odrv12 I__5960 (
            .O(N__27085),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3 ));
    Odrv4 I__5959 (
            .O(N__27082),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3 ));
    CascadeMux I__5958 (
            .O(N__27077),
            .I(N__27074));
    InMux I__5957 (
            .O(N__27074),
            .I(N__27071));
    LocalMux I__5956 (
            .O(N__27071),
            .I(N__27068));
    Odrv12 I__5955 (
            .O(N__27068),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_3 ));
    InMux I__5954 (
            .O(N__27065),
            .I(N__27062));
    LocalMux I__5953 (
            .O(N__27062),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIG6MM1_3 ));
    InMux I__5952 (
            .O(N__27059),
            .I(N__27056));
    LocalMux I__5951 (
            .O(N__27056),
            .I(N__27053));
    Span4Mux_v I__5950 (
            .O(N__27053),
            .I(N__27050));
    Span4Mux_s0_h I__5949 (
            .O(N__27050),
            .I(N__27047));
    Odrv4 I__5948 (
            .O(N__27047),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIASHQ1_2 ));
    CascadeMux I__5947 (
            .O(N__27044),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIC2MM1_2_cascade_ ));
    InMux I__5946 (
            .O(N__27041),
            .I(N__27038));
    LocalMux I__5945 (
            .O(N__27038),
            .I(N__27035));
    Span4Mux_v I__5944 (
            .O(N__27035),
            .I(N__27032));
    Span4Mux_h I__5943 (
            .O(N__27032),
            .I(N__27029));
    Odrv4 I__5942 (
            .O(N__27029),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFHAI8_2 ));
    CascadeMux I__5941 (
            .O(N__27026),
            .I(N__27023));
    InMux I__5940 (
            .O(N__27023),
            .I(N__27020));
    LocalMux I__5939 (
            .O(N__27020),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_2 ));
    InMux I__5938 (
            .O(N__27017),
            .I(N__27014));
    LocalMux I__5937 (
            .O(N__27014),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIS1K32_2 ));
    CascadeMux I__5936 (
            .O(N__27011),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIGEUU1_2_cascade_ ));
    InMux I__5935 (
            .O(N__27008),
            .I(N__27005));
    LocalMux I__5934 (
            .O(N__27005),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_2 ));
    InMux I__5933 (
            .O(N__27002),
            .I(N__26998));
    InMux I__5932 (
            .O(N__27001),
            .I(N__26995));
    LocalMux I__5931 (
            .O(N__26998),
            .I(N__26992));
    LocalMux I__5930 (
            .O(N__26995),
            .I(N__26989));
    Span4Mux_h I__5929 (
            .O(N__26992),
            .I(N__26986));
    Span4Mux_h I__5928 (
            .O(N__26989),
            .I(N__26983));
    Odrv4 I__5927 (
            .O(N__26986),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0 ));
    Odrv4 I__5926 (
            .O(N__26983),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0 ));
    InMux I__5925 (
            .O(N__26978),
            .I(N__26974));
    InMux I__5924 (
            .O(N__26977),
            .I(N__26971));
    LocalMux I__5923 (
            .O(N__26974),
            .I(N__26966));
    LocalMux I__5922 (
            .O(N__26971),
            .I(N__26966));
    Span4Mux_v I__5921 (
            .O(N__26966),
            .I(N__26963));
    Odrv4 I__5920 (
            .O(N__26963),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_1 ));
    InMux I__5919 (
            .O(N__26960),
            .I(N__26957));
    LocalMux I__5918 (
            .O(N__26957),
            .I(N__26953));
    InMux I__5917 (
            .O(N__26956),
            .I(N__26950));
    Odrv4 I__5916 (
            .O(N__26953),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1 ));
    LocalMux I__5915 (
            .O(N__26950),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1 ));
    CascadeMux I__5914 (
            .O(N__26945),
            .I(N__26942));
    InMux I__5913 (
            .O(N__26942),
            .I(N__26939));
    LocalMux I__5912 (
            .O(N__26939),
            .I(N__26936));
    Odrv4 I__5911 (
            .O(N__26936),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_1 ));
    InMux I__5910 (
            .O(N__26933),
            .I(N__26929));
    InMux I__5909 (
            .O(N__26932),
            .I(N__26926));
    LocalMux I__5908 (
            .O(N__26929),
            .I(N__26921));
    LocalMux I__5907 (
            .O(N__26926),
            .I(N__26921));
    Span4Mux_v I__5906 (
            .O(N__26921),
            .I(N__26918));
    Odrv4 I__5905 (
            .O(N__26918),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_2 ));
    InMux I__5904 (
            .O(N__26915),
            .I(N__26911));
    InMux I__5903 (
            .O(N__26914),
            .I(N__26908));
    LocalMux I__5902 (
            .O(N__26911),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2 ));
    LocalMux I__5901 (
            .O(N__26908),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2 ));
    InMux I__5900 (
            .O(N__26903),
            .I(N__26900));
    LocalMux I__5899 (
            .O(N__26900),
            .I(N__26897));
    Span4Mux_h I__5898 (
            .O(N__26897),
            .I(N__26894));
    Odrv4 I__5897 (
            .O(N__26894),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_2 ));
    InMux I__5896 (
            .O(N__26891),
            .I(N__26888));
    LocalMux I__5895 (
            .O(N__26888),
            .I(N__26885));
    IoSpan4Mux I__5894 (
            .O(N__26885),
            .I(N__26882));
    Span4Mux_s3_h I__5893 (
            .O(N__26882),
            .I(N__26878));
    InMux I__5892 (
            .O(N__26881),
            .I(N__26875));
    Sp12to4 I__5891 (
            .O(N__26878),
            .I(N__26870));
    LocalMux I__5890 (
            .O(N__26875),
            .I(N__26870));
    Odrv12 I__5889 (
            .O(N__26870),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_1 ));
    InMux I__5888 (
            .O(N__26867),
            .I(N__26864));
    LocalMux I__5887 (
            .O(N__26864),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_1 ));
    CascadeMux I__5886 (
            .O(N__26861),
            .I(N__26857));
    CascadeMux I__5885 (
            .O(N__26860),
            .I(N__26854));
    InMux I__5884 (
            .O(N__26857),
            .I(N__26851));
    InMux I__5883 (
            .O(N__26854),
            .I(N__26848));
    LocalMux I__5882 (
            .O(N__26851),
            .I(N__26845));
    LocalMux I__5881 (
            .O(N__26848),
            .I(N__26842));
    Span4Mux_v I__5880 (
            .O(N__26845),
            .I(N__26839));
    Span4Mux_v I__5879 (
            .O(N__26842),
            .I(N__26836));
    Span4Mux_v I__5878 (
            .O(N__26839),
            .I(N__26833));
    Span4Mux_h I__5877 (
            .O(N__26836),
            .I(N__26830));
    Odrv4 I__5876 (
            .O(N__26833),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1 ));
    Odrv4 I__5875 (
            .O(N__26830),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1 ));
    InMux I__5874 (
            .O(N__26825),
            .I(N__26822));
    LocalMux I__5873 (
            .O(N__26822),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_295 ));
    InMux I__5872 (
            .O(N__26819),
            .I(N__26816));
    LocalMux I__5871 (
            .O(N__26816),
            .I(N__26813));
    Span4Mux_v I__5870 (
            .O(N__26813),
            .I(N__26809));
    InMux I__5869 (
            .O(N__26812),
            .I(N__26806));
    Odrv4 I__5868 (
            .O(N__26809),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1 ));
    LocalMux I__5867 (
            .O(N__26806),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1 ));
    CascadeMux I__5866 (
            .O(N__26801),
            .I(N__26798));
    InMux I__5865 (
            .O(N__26798),
            .I(N__26795));
    LocalMux I__5864 (
            .O(N__26795),
            .I(N__26791));
    InMux I__5863 (
            .O(N__26794),
            .I(N__26788));
    Odrv4 I__5862 (
            .O(N__26791),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1 ));
    LocalMux I__5861 (
            .O(N__26788),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1 ));
    CascadeMux I__5860 (
            .O(N__26783),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_1_cascade_ ));
    InMux I__5859 (
            .O(N__26780),
            .I(N__26777));
    LocalMux I__5858 (
            .O(N__26777),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_215 ));
    InMux I__5857 (
            .O(N__26774),
            .I(N__26771));
    LocalMux I__5856 (
            .O(N__26771),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_1 ));
    CascadeMux I__5855 (
            .O(N__26768),
            .I(N__26765));
    InMux I__5854 (
            .O(N__26765),
            .I(N__26762));
    LocalMux I__5853 (
            .O(N__26762),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_239 ));
    CascadeMux I__5852 (
            .O(N__26759),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_2_cascade_ ));
    InMux I__5851 (
            .O(N__26756),
            .I(N__26753));
    LocalMux I__5850 (
            .O(N__26753),
            .I(N__26749));
    InMux I__5849 (
            .O(N__26752),
            .I(N__26746));
    Odrv4 I__5848 (
            .O(N__26749),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2 ));
    LocalMux I__5847 (
            .O(N__26746),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2 ));
    CascadeMux I__5846 (
            .O(N__26741),
            .I(N__26738));
    InMux I__5845 (
            .O(N__26738),
            .I(N__26735));
    LocalMux I__5844 (
            .O(N__26735),
            .I(N__26732));
    Span4Mux_s2_h I__5843 (
            .O(N__26732),
            .I(N__26728));
    InMux I__5842 (
            .O(N__26731),
            .I(N__26725));
    Odrv4 I__5841 (
            .O(N__26728),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2 ));
    LocalMux I__5840 (
            .O(N__26725),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2 ));
    InMux I__5839 (
            .O(N__26720),
            .I(N__26717));
    LocalMux I__5838 (
            .O(N__26717),
            .I(N__26713));
    InMux I__5837 (
            .O(N__26716),
            .I(N__26710));
    Odrv4 I__5836 (
            .O(N__26713),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2 ));
    LocalMux I__5835 (
            .O(N__26710),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2 ));
    CascadeMux I__5834 (
            .O(N__26705),
            .I(N__26702));
    InMux I__5833 (
            .O(N__26702),
            .I(N__26699));
    LocalMux I__5832 (
            .O(N__26699),
            .I(N__26696));
    Span4Mux_v I__5831 (
            .O(N__26696),
            .I(N__26693));
    Odrv4 I__5830 (
            .O(N__26693),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_2 ));
    InMux I__5829 (
            .O(N__26690),
            .I(N__26686));
    InMux I__5828 (
            .O(N__26689),
            .I(N__26683));
    LocalMux I__5827 (
            .O(N__26686),
            .I(N__26680));
    LocalMux I__5826 (
            .O(N__26683),
            .I(N__26677));
    Span4Mux_h I__5825 (
            .O(N__26680),
            .I(N__26674));
    Odrv12 I__5824 (
            .O(N__26677),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4 ));
    Odrv4 I__5823 (
            .O(N__26674),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4 ));
    CascadeMux I__5822 (
            .O(N__26669),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_4_cascade_ ));
    InMux I__5821 (
            .O(N__26666),
            .I(N__26663));
    LocalMux I__5820 (
            .O(N__26663),
            .I(N__26660));
    Span4Mux_v I__5819 (
            .O(N__26660),
            .I(N__26657));
    Span4Mux_h I__5818 (
            .O(N__26657),
            .I(N__26654));
    Odrv4 I__5817 (
            .O(N__26654),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIKAMM1_4 ));
    CascadeMux I__5816 (
            .O(N__26651),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_1_cascade_ ));
    InMux I__5815 (
            .O(N__26648),
            .I(N__26644));
    InMux I__5814 (
            .O(N__26647),
            .I(N__26641));
    LocalMux I__5813 (
            .O(N__26644),
            .I(N__26638));
    LocalMux I__5812 (
            .O(N__26641),
            .I(N__26635));
    Span4Mux_v I__5811 (
            .O(N__26638),
            .I(N__26632));
    Span12Mux_s3_h I__5810 (
            .O(N__26635),
            .I(N__26629));
    Odrv4 I__5809 (
            .O(N__26632),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2 ));
    Odrv12 I__5808 (
            .O(N__26629),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2 ));
    CascadeMux I__5807 (
            .O(N__26624),
            .I(N__26621));
    InMux I__5806 (
            .O(N__26621),
            .I(N__26617));
    InMux I__5805 (
            .O(N__26620),
            .I(N__26614));
    LocalMux I__5804 (
            .O(N__26617),
            .I(N__26609));
    LocalMux I__5803 (
            .O(N__26614),
            .I(N__26609));
    Odrv12 I__5802 (
            .O(N__26609),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_2 ));
    CascadeMux I__5801 (
            .O(N__26606),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_2_cascade_ ));
    InMux I__5800 (
            .O(N__26603),
            .I(N__26599));
    InMux I__5799 (
            .O(N__26602),
            .I(N__26596));
    LocalMux I__5798 (
            .O(N__26599),
            .I(N__26593));
    LocalMux I__5797 (
            .O(N__26596),
            .I(N__26590));
    Span4Mux_s2_h I__5796 (
            .O(N__26593),
            .I(N__26587));
    Span4Mux_s2_h I__5795 (
            .O(N__26590),
            .I(N__26584));
    Odrv4 I__5794 (
            .O(N__26587),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2 ));
    Odrv4 I__5793 (
            .O(N__26584),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2 ));
    InMux I__5792 (
            .O(N__26579),
            .I(N__26575));
    InMux I__5791 (
            .O(N__26578),
            .I(N__26572));
    LocalMux I__5790 (
            .O(N__26575),
            .I(N__26569));
    LocalMux I__5789 (
            .O(N__26572),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1 ));
    Odrv12 I__5788 (
            .O(N__26569),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1 ));
    CascadeMux I__5787 (
            .O(N__26564),
            .I(N__26561));
    InMux I__5786 (
            .O(N__26561),
            .I(N__26558));
    LocalMux I__5785 (
            .O(N__26558),
            .I(N__26555));
    Odrv12 I__5784 (
            .O(N__26555),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_1 ));
    InMux I__5783 (
            .O(N__26552),
            .I(N__26549));
    LocalMux I__5782 (
            .O(N__26549),
            .I(N__26546));
    Span4Mux_h I__5781 (
            .O(N__26546),
            .I(N__26543));
    Odrv4 I__5780 (
            .O(N__26543),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1 ));
    InMux I__5779 (
            .O(N__26540),
            .I(N__26537));
    LocalMux I__5778 (
            .O(N__26537),
            .I(N__26533));
    InMux I__5777 (
            .O(N__26536),
            .I(N__26530));
    Span4Mux_v I__5776 (
            .O(N__26533),
            .I(N__26527));
    LocalMux I__5775 (
            .O(N__26530),
            .I(N__26524));
    Odrv4 I__5774 (
            .O(N__26527),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1 ));
    Odrv12 I__5773 (
            .O(N__26524),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1 ));
    CascadeMux I__5772 (
            .O(N__26519),
            .I(N__26516));
    InMux I__5771 (
            .O(N__26516),
            .I(N__26512));
    CascadeMux I__5770 (
            .O(N__26515),
            .I(N__26509));
    LocalMux I__5769 (
            .O(N__26512),
            .I(N__26506));
    InMux I__5768 (
            .O(N__26509),
            .I(N__26503));
    Span4Mux_v I__5767 (
            .O(N__26506),
            .I(N__26500));
    LocalMux I__5766 (
            .O(N__26503),
            .I(N__26497));
    Span4Mux_v I__5765 (
            .O(N__26500),
            .I(N__26494));
    Odrv12 I__5764 (
            .O(N__26497),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1 ));
    Odrv4 I__5763 (
            .O(N__26494),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1 ));
    InMux I__5762 (
            .O(N__26489),
            .I(N__26486));
    LocalMux I__5761 (
            .O(N__26486),
            .I(N__26483));
    Odrv12 I__5760 (
            .O(N__26483),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_271 ));
    CascadeMux I__5759 (
            .O(N__26480),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_1_cascade_ ));
    InMux I__5758 (
            .O(N__26477),
            .I(N__26474));
    LocalMux I__5757 (
            .O(N__26474),
            .I(N__26471));
    Span4Mux_h I__5756 (
            .O(N__26471),
            .I(N__26468));
    Span4Mux_h I__5755 (
            .O(N__26468),
            .I(N__26465));
    Odrv4 I__5754 (
            .O(N__26465),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_311 ));
    InMux I__5753 (
            .O(N__26462),
            .I(N__26459));
    LocalMux I__5752 (
            .O(N__26459),
            .I(N__26455));
    InMux I__5751 (
            .O(N__26458),
            .I(N__26452));
    Span4Mux_v I__5750 (
            .O(N__26455),
            .I(N__26447));
    LocalMux I__5749 (
            .O(N__26452),
            .I(N__26447));
    Odrv4 I__5748 (
            .O(N__26447),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_0 ));
    InMux I__5747 (
            .O(N__26444),
            .I(N__26440));
    InMux I__5746 (
            .O(N__26443),
            .I(N__26437));
    LocalMux I__5745 (
            .O(N__26440),
            .I(N__26434));
    LocalMux I__5744 (
            .O(N__26437),
            .I(N__26431));
    Span4Mux_h I__5743 (
            .O(N__26434),
            .I(N__26428));
    Span4Mux_h I__5742 (
            .O(N__26431),
            .I(N__26425));
    Odrv4 I__5741 (
            .O(N__26428),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5 ));
    Odrv4 I__5740 (
            .O(N__26425),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5 ));
    InMux I__5739 (
            .O(N__26420),
            .I(N__26414));
    InMux I__5738 (
            .O(N__26419),
            .I(N__26414));
    LocalMux I__5737 (
            .O(N__26414),
            .I(N__26411));
    Span12Mux_s6_v I__5736 (
            .O(N__26411),
            .I(N__26408));
    Odrv12 I__5735 (
            .O(N__26408),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_6 ));
    CEMux I__5734 (
            .O(N__26405),
            .I(N__26402));
    LocalMux I__5733 (
            .O(N__26402),
            .I(N__26399));
    Span4Mux_v I__5732 (
            .O(N__26399),
            .I(N__26396));
    Span4Mux_h I__5731 (
            .O(N__26396),
            .I(N__26393));
    Odrv4 I__5730 (
            .O(N__26393),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe27 ));
    InMux I__5729 (
            .O(N__26390),
            .I(N__26387));
    LocalMux I__5728 (
            .O(N__26387),
            .I(N__26384));
    Span4Mux_s3_h I__5727 (
            .O(N__26384),
            .I(N__26380));
    InMux I__5726 (
            .O(N__26383),
            .I(N__26377));
    Odrv4 I__5725 (
            .O(N__26380),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3 ));
    LocalMux I__5724 (
            .O(N__26377),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3 ));
    CascadeMux I__5723 (
            .O(N__26372),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_3_cascade_ ));
    InMux I__5722 (
            .O(N__26369),
            .I(N__26366));
    LocalMux I__5721 (
            .O(N__26366),
            .I(N__26362));
    InMux I__5720 (
            .O(N__26365),
            .I(N__26359));
    Odrv4 I__5719 (
            .O(N__26362),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3 ));
    LocalMux I__5718 (
            .O(N__26359),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3 ));
    CascadeMux I__5717 (
            .O(N__26354),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_2_cascade_ ));
    InMux I__5716 (
            .O(N__26351),
            .I(N__26348));
    LocalMux I__5715 (
            .O(N__26348),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_2 ));
    CascadeMux I__5714 (
            .O(N__26345),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_2_cascade_ ));
    InMux I__5713 (
            .O(N__26342),
            .I(N__26339));
    LocalMux I__5712 (
            .O(N__26339),
            .I(N__26336));
    Span4Mux_h I__5711 (
            .O(N__26336),
            .I(N__26333));
    Span4Mux_v I__5710 (
            .O(N__26333),
            .I(N__26330));
    Odrv4 I__5709 (
            .O(N__26330),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_2 ));
    InMux I__5708 (
            .O(N__26327),
            .I(N__26324));
    LocalMux I__5707 (
            .O(N__26324),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_2 ));
    InMux I__5706 (
            .O(N__26321),
            .I(N__26318));
    LocalMux I__5705 (
            .O(N__26318),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_2 ));
    InMux I__5704 (
            .O(N__26315),
            .I(N__26311));
    InMux I__5703 (
            .O(N__26314),
            .I(N__26308));
    LocalMux I__5702 (
            .O(N__26311),
            .I(N__26305));
    LocalMux I__5701 (
            .O(N__26308),
            .I(N__26302));
    Span4Mux_h I__5700 (
            .O(N__26305),
            .I(N__26297));
    Span4Mux_h I__5699 (
            .O(N__26302),
            .I(N__26297));
    Odrv4 I__5698 (
            .O(N__26297),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_6 ));
    CEMux I__5697 (
            .O(N__26294),
            .I(N__26291));
    LocalMux I__5696 (
            .O(N__26291),
            .I(N__26288));
    Sp12to4 I__5695 (
            .O(N__26288),
            .I(N__26285));
    Odrv12 I__5694 (
            .O(N__26285),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe29 ));
    CascadeMux I__5693 (
            .O(N__26282),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_3_cascade_ ));
    InMux I__5692 (
            .O(N__26279),
            .I(N__26276));
    LocalMux I__5691 (
            .O(N__26276),
            .I(N__26273));
    Odrv4 I__5690 (
            .O(N__26273),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_3 ));
    CascadeMux I__5689 (
            .O(N__26270),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_3_cascade_ ));
    CascadeMux I__5688 (
            .O(N__26267),
            .I(N__26264));
    InMux I__5687 (
            .O(N__26264),
            .I(N__26261));
    LocalMux I__5686 (
            .O(N__26261),
            .I(N__26258));
    Span4Mux_h I__5685 (
            .O(N__26258),
            .I(N__26255));
    Span4Mux_v I__5684 (
            .O(N__26255),
            .I(N__26252));
    Span4Mux_v I__5683 (
            .O(N__26252),
            .I(N__26249));
    Odrv4 I__5682 (
            .O(N__26249),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_3 ));
    InMux I__5681 (
            .O(N__26246),
            .I(N__26243));
    LocalMux I__5680 (
            .O(N__26243),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_3 ));
    InMux I__5679 (
            .O(N__26240),
            .I(N__26237));
    LocalMux I__5678 (
            .O(N__26237),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_3 ));
    InMux I__5677 (
            .O(N__26234),
            .I(N__26228));
    InMux I__5676 (
            .O(N__26233),
            .I(N__26228));
    LocalMux I__5675 (
            .O(N__26228),
            .I(N__26225));
    Span4Mux_s2_h I__5674 (
            .O(N__26225),
            .I(N__26222));
    Odrv4 I__5673 (
            .O(N__26222),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_3 ));
    CascadeMux I__5672 (
            .O(N__26219),
            .I(N__26216));
    InMux I__5671 (
            .O(N__26216),
            .I(N__26210));
    InMux I__5670 (
            .O(N__26215),
            .I(N__26210));
    LocalMux I__5669 (
            .O(N__26210),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_3 ));
    InMux I__5668 (
            .O(N__26207),
            .I(N__26204));
    LocalMux I__5667 (
            .O(N__26204),
            .I(N__26201));
    Span4Mux_h I__5666 (
            .O(N__26201),
            .I(N__26197));
    InMux I__5665 (
            .O(N__26200),
            .I(N__26194));
    Odrv4 I__5664 (
            .O(N__26197),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3 ));
    LocalMux I__5663 (
            .O(N__26194),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3 ));
    InMux I__5662 (
            .O(N__26189),
            .I(N__26186));
    LocalMux I__5661 (
            .O(N__26186),
            .I(N__26182));
    InMux I__5660 (
            .O(N__26185),
            .I(N__26179));
    Span4Mux_v I__5659 (
            .O(N__26182),
            .I(N__26176));
    LocalMux I__5658 (
            .O(N__26179),
            .I(N__26173));
    Odrv4 I__5657 (
            .O(N__26176),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4 ));
    Odrv4 I__5656 (
            .O(N__26173),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4 ));
    CEMux I__5655 (
            .O(N__26168),
            .I(N__26164));
    CEMux I__5654 (
            .O(N__26167),
            .I(N__26161));
    LocalMux I__5653 (
            .O(N__26164),
            .I(N__26157));
    LocalMux I__5652 (
            .O(N__26161),
            .I(N__26154));
    CEMux I__5651 (
            .O(N__26160),
            .I(N__26151));
    Sp12to4 I__5650 (
            .O(N__26157),
            .I(N__26148));
    Span4Mux_s3_v I__5649 (
            .O(N__26154),
            .I(N__26145));
    LocalMux I__5648 (
            .O(N__26151),
            .I(N__26142));
    Span12Mux_s5_h I__5647 (
            .O(N__26148),
            .I(N__26139));
    Span4Mux_h I__5646 (
            .O(N__26145),
            .I(N__26136));
    Span4Mux_h I__5645 (
            .O(N__26142),
            .I(N__26133));
    Odrv12 I__5644 (
            .O(N__26139),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3 ));
    Odrv4 I__5643 (
            .O(N__26136),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3 ));
    Odrv4 I__5642 (
            .O(N__26133),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3 ));
    InMux I__5641 (
            .O(N__26126),
            .I(N__26122));
    InMux I__5640 (
            .O(N__26125),
            .I(N__26119));
    LocalMux I__5639 (
            .O(N__26122),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5 ));
    LocalMux I__5638 (
            .O(N__26119),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5 ));
    InMux I__5637 (
            .O(N__26114),
            .I(N__26110));
    InMux I__5636 (
            .O(N__26113),
            .I(N__26107));
    LocalMux I__5635 (
            .O(N__26110),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5 ));
    LocalMux I__5634 (
            .O(N__26107),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5 ));
    InMux I__5633 (
            .O(N__26102),
            .I(N__26099));
    LocalMux I__5632 (
            .O(N__26099),
            .I(N__26096));
    Span4Mux_v I__5631 (
            .O(N__26096),
            .I(N__26093));
    Odrv4 I__5630 (
            .O(N__26093),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_5 ));
    InMux I__5629 (
            .O(N__26090),
            .I(N__26084));
    InMux I__5628 (
            .O(N__26089),
            .I(N__26084));
    LocalMux I__5627 (
            .O(N__26084),
            .I(N__26081));
    Span4Mux_v I__5626 (
            .O(N__26081),
            .I(N__26078));
    Odrv4 I__5625 (
            .O(N__26078),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_0 ));
    InMux I__5624 (
            .O(N__26075),
            .I(N__26071));
    CascadeMux I__5623 (
            .O(N__26074),
            .I(N__26068));
    LocalMux I__5622 (
            .O(N__26071),
            .I(N__26065));
    InMux I__5621 (
            .O(N__26068),
            .I(N__26062));
    Span4Mux_v I__5620 (
            .O(N__26065),
            .I(N__26057));
    LocalMux I__5619 (
            .O(N__26062),
            .I(N__26057));
    Span4Mux_h I__5618 (
            .O(N__26057),
            .I(N__26054));
    Odrv4 I__5617 (
            .O(N__26054),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_4 ));
    InMux I__5616 (
            .O(N__26051),
            .I(N__26045));
    InMux I__5615 (
            .O(N__26050),
            .I(N__26045));
    LocalMux I__5614 (
            .O(N__26045),
            .I(N__26042));
    Span4Mux_v I__5613 (
            .O(N__26042),
            .I(N__26039));
    Span4Mux_h I__5612 (
            .O(N__26039),
            .I(N__26036));
    Odrv4 I__5611 (
            .O(N__26036),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_5 ));
    InMux I__5610 (
            .O(N__26033),
            .I(N__26029));
    InMux I__5609 (
            .O(N__26032),
            .I(N__26026));
    LocalMux I__5608 (
            .O(N__26029),
            .I(N__26023));
    LocalMux I__5607 (
            .O(N__26026),
            .I(N__26020));
    Span4Mux_h I__5606 (
            .O(N__26023),
            .I(N__26017));
    Span4Mux_h I__5605 (
            .O(N__26020),
            .I(N__26014));
    Odrv4 I__5604 (
            .O(N__26017),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1 ));
    Odrv4 I__5603 (
            .O(N__26014),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1 ));
    InMux I__5602 (
            .O(N__26009),
            .I(N__26006));
    LocalMux I__5601 (
            .O(N__26006),
            .I(N__26003));
    Span4Mux_h I__5600 (
            .O(N__26003),
            .I(N__25999));
    InMux I__5599 (
            .O(N__26002),
            .I(N__25996));
    Odrv4 I__5598 (
            .O(N__25999),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2 ));
    LocalMux I__5597 (
            .O(N__25996),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2 ));
    InMux I__5596 (
            .O(N__25991),
            .I(N__25988));
    LocalMux I__5595 (
            .O(N__25988),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_2 ));
    InMux I__5594 (
            .O(N__25985),
            .I(N__25982));
    LocalMux I__5593 (
            .O(N__25982),
            .I(N__25978));
    InMux I__5592 (
            .O(N__25981),
            .I(N__25975));
    Odrv4 I__5591 (
            .O(N__25978),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3 ));
    LocalMux I__5590 (
            .O(N__25975),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3 ));
    InMux I__5589 (
            .O(N__25970),
            .I(N__25967));
    LocalMux I__5588 (
            .O(N__25967),
            .I(N__25964));
    Span4Mux_h I__5587 (
            .O(N__25964),
            .I(N__25961));
    Odrv4 I__5586 (
            .O(N__25961),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_3 ));
    CEMux I__5585 (
            .O(N__25958),
            .I(N__25954));
    CEMux I__5584 (
            .O(N__25957),
            .I(N__25951));
    LocalMux I__5583 (
            .O(N__25954),
            .I(N__25948));
    LocalMux I__5582 (
            .O(N__25951),
            .I(N__25945));
    Span4Mux_v I__5581 (
            .O(N__25948),
            .I(N__25941));
    Span4Mux_s3_v I__5580 (
            .O(N__25945),
            .I(N__25938));
    CEMux I__5579 (
            .O(N__25944),
            .I(N__25935));
    Span4Mux_h I__5578 (
            .O(N__25941),
            .I(N__25932));
    Sp12to4 I__5577 (
            .O(N__25938),
            .I(N__25929));
    LocalMux I__5576 (
            .O(N__25935),
            .I(N__25926));
    Sp12to4 I__5575 (
            .O(N__25932),
            .I(N__25921));
    Span12Mux_s8_h I__5574 (
            .O(N__25929),
            .I(N__25921));
    Span4Mux_v I__5573 (
            .O(N__25926),
            .I(N__25918));
    Odrv12 I__5572 (
            .O(N__25921),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2 ));
    Odrv4 I__5571 (
            .O(N__25918),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2 ));
    InMux I__5570 (
            .O(N__25913),
            .I(N__25909));
    InMux I__5569 (
            .O(N__25912),
            .I(N__25906));
    LocalMux I__5568 (
            .O(N__25909),
            .I(N__25903));
    LocalMux I__5567 (
            .O(N__25906),
            .I(N__25900));
    Span4Mux_h I__5566 (
            .O(N__25903),
            .I(N__25897));
    Span4Mux_h I__5565 (
            .O(N__25900),
            .I(N__25894));
    Span4Mux_v I__5564 (
            .O(N__25897),
            .I(N__25891));
    Span4Mux_v I__5563 (
            .O(N__25894),
            .I(N__25888));
    Odrv4 I__5562 (
            .O(N__25891),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0 ));
    Odrv4 I__5561 (
            .O(N__25888),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0 ));
    InMux I__5560 (
            .O(N__25883),
            .I(N__25879));
    InMux I__5559 (
            .O(N__25882),
            .I(N__25876));
    LocalMux I__5558 (
            .O(N__25879),
            .I(N__25873));
    LocalMux I__5557 (
            .O(N__25876),
            .I(N__25870));
    Span4Mux_h I__5556 (
            .O(N__25873),
            .I(N__25867));
    Span4Mux_v I__5555 (
            .O(N__25870),
            .I(N__25864));
    Odrv4 I__5554 (
            .O(N__25867),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1 ));
    Odrv4 I__5553 (
            .O(N__25864),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1 ));
    InMux I__5552 (
            .O(N__25859),
            .I(N__25856));
    LocalMux I__5551 (
            .O(N__25856),
            .I(N__25853));
    Span4Mux_v I__5550 (
            .O(N__25853),
            .I(N__25850));
    Span4Mux_s1_v I__5549 (
            .O(N__25850),
            .I(N__25846));
    InMux I__5548 (
            .O(N__25849),
            .I(N__25843));
    Odrv4 I__5547 (
            .O(N__25846),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2 ));
    LocalMux I__5546 (
            .O(N__25843),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2 ));
    InMux I__5545 (
            .O(N__25838),
            .I(N__25835));
    LocalMux I__5544 (
            .O(N__25835),
            .I(N__25832));
    Odrv4 I__5543 (
            .O(N__25832),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_2 ));
    CascadeMux I__5542 (
            .O(N__25829),
            .I(N__25826));
    InMux I__5541 (
            .O(N__25826),
            .I(N__25823));
    LocalMux I__5540 (
            .O(N__25823),
            .I(N__25820));
    Span4Mux_v I__5539 (
            .O(N__25820),
            .I(N__25817));
    Odrv4 I__5538 (
            .O(N__25817),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_2 ));
    InMux I__5537 (
            .O(N__25814),
            .I(N__25811));
    LocalMux I__5536 (
            .O(N__25811),
            .I(N__25808));
    Span4Mux_v I__5535 (
            .O(N__25808),
            .I(N__25805));
    Span4Mux_h I__5534 (
            .O(N__25805),
            .I(N__25802));
    Odrv4 I__5533 (
            .O(N__25802),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_2 ));
    CascadeMux I__5532 (
            .O(N__25799),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_2_cascade_ ));
    SRMux I__5531 (
            .O(N__25796),
            .I(N__25793));
    LocalMux I__5530 (
            .O(N__25793),
            .I(N__25789));
    InMux I__5529 (
            .O(N__25792),
            .I(N__25786));
    Span4Mux_h I__5528 (
            .O(N__25789),
            .I(N__25777));
    LocalMux I__5527 (
            .O(N__25786),
            .I(N__25777));
    InMux I__5526 (
            .O(N__25785),
            .I(N__25774));
    InMux I__5525 (
            .O(N__25784),
            .I(N__25770));
    InMux I__5524 (
            .O(N__25783),
            .I(N__25767));
    InMux I__5523 (
            .O(N__25782),
            .I(N__25764));
    Span4Mux_v I__5522 (
            .O(N__25777),
            .I(N__25756));
    LocalMux I__5521 (
            .O(N__25774),
            .I(N__25756));
    InMux I__5520 (
            .O(N__25773),
            .I(N__25752));
    LocalMux I__5519 (
            .O(N__25770),
            .I(N__25749));
    LocalMux I__5518 (
            .O(N__25767),
            .I(N__25744));
    LocalMux I__5517 (
            .O(N__25764),
            .I(N__25744));
    InMux I__5516 (
            .O(N__25763),
            .I(N__25741));
    InMux I__5515 (
            .O(N__25762),
            .I(N__25738));
    InMux I__5514 (
            .O(N__25761),
            .I(N__25734));
    Span4Mux_h I__5513 (
            .O(N__25756),
            .I(N__25731));
    InMux I__5512 (
            .O(N__25755),
            .I(N__25728));
    LocalMux I__5511 (
            .O(N__25752),
            .I(N__25725));
    Span4Mux_v I__5510 (
            .O(N__25749),
            .I(N__25720));
    Span4Mux_v I__5509 (
            .O(N__25744),
            .I(N__25720));
    LocalMux I__5508 (
            .O(N__25741),
            .I(N__25715));
    LocalMux I__5507 (
            .O(N__25738),
            .I(N__25715));
    InMux I__5506 (
            .O(N__25737),
            .I(N__25712));
    LocalMux I__5505 (
            .O(N__25734),
            .I(N__25709));
    Span4Mux_v I__5504 (
            .O(N__25731),
            .I(N__25706));
    LocalMux I__5503 (
            .O(N__25728),
            .I(N__25703));
    Span4Mux_v I__5502 (
            .O(N__25725),
            .I(N__25700));
    Span4Mux_h I__5501 (
            .O(N__25720),
            .I(N__25693));
    Span4Mux_v I__5500 (
            .O(N__25715),
            .I(N__25693));
    LocalMux I__5499 (
            .O(N__25712),
            .I(N__25693));
    Span12Mux_s9_h I__5498 (
            .O(N__25709),
            .I(N__25690));
    Span4Mux_h I__5497 (
            .O(N__25706),
            .I(N__25685));
    Span4Mux_v I__5496 (
            .O(N__25703),
            .I(N__25685));
    Span4Mux_s2_h I__5495 (
            .O(N__25700),
            .I(N__25680));
    Span4Mux_h I__5494 (
            .O(N__25693),
            .I(N__25680));
    Odrv12 I__5493 (
            .O(N__25690),
            .I(instruction_7));
    Odrv4 I__5492 (
            .O(N__25685),
            .I(instruction_7));
    Odrv4 I__5491 (
            .O(N__25680),
            .I(instruction_7));
    CascadeMux I__5490 (
            .O(N__25673),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_2_cascade_ ));
    InMux I__5489 (
            .O(N__25670),
            .I(N__25662));
    InMux I__5488 (
            .O(N__25669),
            .I(N__25662));
    InMux I__5487 (
            .O(N__25668),
            .I(N__25653));
    InMux I__5486 (
            .O(N__25667),
            .I(N__25653));
    LocalMux I__5485 (
            .O(N__25662),
            .I(N__25650));
    InMux I__5484 (
            .O(N__25661),
            .I(N__25645));
    InMux I__5483 (
            .O(N__25660),
            .I(N__25645));
    InMux I__5482 (
            .O(N__25659),
            .I(N__25640));
    InMux I__5481 (
            .O(N__25658),
            .I(N__25640));
    LocalMux I__5480 (
            .O(N__25653),
            .I(N__25632));
    Span4Mux_h I__5479 (
            .O(N__25650),
            .I(N__25627));
    LocalMux I__5478 (
            .O(N__25645),
            .I(N__25627));
    LocalMux I__5477 (
            .O(N__25640),
            .I(N__25624));
    InMux I__5476 (
            .O(N__25639),
            .I(N__25619));
    InMux I__5475 (
            .O(N__25638),
            .I(N__25619));
    InMux I__5474 (
            .O(N__25637),
            .I(N__25616));
    InMux I__5473 (
            .O(N__25636),
            .I(N__25613));
    InMux I__5472 (
            .O(N__25635),
            .I(N__25610));
    Span4Mux_h I__5471 (
            .O(N__25632),
            .I(N__25606));
    Span4Mux_v I__5470 (
            .O(N__25627),
            .I(N__25598));
    Span4Mux_v I__5469 (
            .O(N__25624),
            .I(N__25593));
    LocalMux I__5468 (
            .O(N__25619),
            .I(N__25593));
    LocalMux I__5467 (
            .O(N__25616),
            .I(N__25590));
    LocalMux I__5466 (
            .O(N__25613),
            .I(N__25585));
    LocalMux I__5465 (
            .O(N__25610),
            .I(N__25585));
    InMux I__5464 (
            .O(N__25609),
            .I(N__25582));
    Span4Mux_v I__5463 (
            .O(N__25606),
            .I(N__25579));
    InMux I__5462 (
            .O(N__25605),
            .I(N__25574));
    InMux I__5461 (
            .O(N__25604),
            .I(N__25574));
    InMux I__5460 (
            .O(N__25603),
            .I(N__25571));
    InMux I__5459 (
            .O(N__25602),
            .I(N__25566));
    InMux I__5458 (
            .O(N__25601),
            .I(N__25566));
    Span4Mux_h I__5457 (
            .O(N__25598),
            .I(N__25561));
    Span4Mux_h I__5456 (
            .O(N__25593),
            .I(N__25561));
    Span4Mux_h I__5455 (
            .O(N__25590),
            .I(N__25556));
    Span4Mux_h I__5454 (
            .O(N__25585),
            .I(N__25556));
    LocalMux I__5453 (
            .O(N__25582),
            .I(\processor_zipi8.bank ));
    Odrv4 I__5452 (
            .O(N__25579),
            .I(\processor_zipi8.bank ));
    LocalMux I__5451 (
            .O(N__25574),
            .I(\processor_zipi8.bank ));
    LocalMux I__5450 (
            .O(N__25571),
            .I(\processor_zipi8.bank ));
    LocalMux I__5449 (
            .O(N__25566),
            .I(\processor_zipi8.bank ));
    Odrv4 I__5448 (
            .O(N__25561),
            .I(\processor_zipi8.bank ));
    Odrv4 I__5447 (
            .O(N__25556),
            .I(\processor_zipi8.bank ));
    InMux I__5446 (
            .O(N__25541),
            .I(N__25537));
    CascadeMux I__5445 (
            .O(N__25540),
            .I(N__25534));
    LocalMux I__5444 (
            .O(N__25537),
            .I(N__25531));
    InMux I__5443 (
            .O(N__25534),
            .I(N__25528));
    Span4Mux_v I__5442 (
            .O(N__25531),
            .I(N__25525));
    LocalMux I__5441 (
            .O(N__25528),
            .I(N__25522));
    Span4Mux_v I__5440 (
            .O(N__25525),
            .I(N__25517));
    Span4Mux_s3_h I__5439 (
            .O(N__25522),
            .I(N__25517));
    Span4Mux_s3_v I__5438 (
            .O(N__25517),
            .I(N__25514));
    Span4Mux_h I__5437 (
            .O(N__25514),
            .I(N__25511));
    Odrv4 I__5436 (
            .O(N__25511),
            .I(\processor_zipi8.sy_2 ));
    CascadeMux I__5435 (
            .O(N__25508),
            .I(N__25505));
    InMux I__5434 (
            .O(N__25505),
            .I(N__25501));
    InMux I__5433 (
            .O(N__25504),
            .I(N__25498));
    LocalMux I__5432 (
            .O(N__25501),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2 ));
    LocalMux I__5431 (
            .O(N__25498),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2 ));
    InMux I__5430 (
            .O(N__25493),
            .I(N__25490));
    LocalMux I__5429 (
            .O(N__25490),
            .I(N__25486));
    InMux I__5428 (
            .O(N__25489),
            .I(N__25483));
    Span4Mux_h I__5427 (
            .O(N__25486),
            .I(N__25480));
    LocalMux I__5426 (
            .O(N__25483),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2 ));
    Odrv4 I__5425 (
            .O(N__25480),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2 ));
    CascadeMux I__5424 (
            .O(N__25475),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_2_cascade_ ));
    InMux I__5423 (
            .O(N__25472),
            .I(N__25469));
    LocalMux I__5422 (
            .O(N__25469),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_2 ));
    InMux I__5421 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__5420 (
            .O(N__25463),
            .I(N__25460));
    Odrv4 I__5419 (
            .O(N__25460),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_2 ));
    CascadeMux I__5418 (
            .O(N__25457),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_2_cascade_ ));
    InMux I__5417 (
            .O(N__25454),
            .I(N__25451));
    LocalMux I__5416 (
            .O(N__25451),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_2 ));
    InMux I__5415 (
            .O(N__25448),
            .I(N__25444));
    InMux I__5414 (
            .O(N__25447),
            .I(N__25441));
    LocalMux I__5413 (
            .O(N__25444),
            .I(N__25438));
    LocalMux I__5412 (
            .O(N__25441),
            .I(N__25435));
    Span4Mux_v I__5411 (
            .O(N__25438),
            .I(N__25430));
    Span4Mux_v I__5410 (
            .O(N__25435),
            .I(N__25430));
    Span4Mux_v I__5409 (
            .O(N__25430),
            .I(N__25427));
    Odrv4 I__5408 (
            .O(N__25427),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_0 ));
    InMux I__5407 (
            .O(N__25424),
            .I(N__25420));
    InMux I__5406 (
            .O(N__25423),
            .I(N__25417));
    LocalMux I__5405 (
            .O(N__25420),
            .I(N__25414));
    LocalMux I__5404 (
            .O(N__25417),
            .I(N__25411));
    Odrv4 I__5403 (
            .O(N__25414),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1 ));
    Odrv4 I__5402 (
            .O(N__25411),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1 ));
    CascadeMux I__5401 (
            .O(N__25406),
            .I(N__25402));
    InMux I__5400 (
            .O(N__25405),
            .I(N__25399));
    InMux I__5399 (
            .O(N__25402),
            .I(N__25396));
    LocalMux I__5398 (
            .O(N__25399),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1 ));
    LocalMux I__5397 (
            .O(N__25396),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1 ));
    InMux I__5396 (
            .O(N__25391),
            .I(N__25387));
    InMux I__5395 (
            .O(N__25390),
            .I(N__25384));
    LocalMux I__5394 (
            .O(N__25387),
            .I(N__25379));
    LocalMux I__5393 (
            .O(N__25384),
            .I(N__25379));
    Span4Mux_h I__5392 (
            .O(N__25379),
            .I(N__25376));
    Odrv4 I__5391 (
            .O(N__25376),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_1 ));
    CascadeMux I__5390 (
            .O(N__25373),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_1_cascade_ ));
    InMux I__5389 (
            .O(N__25370),
            .I(N__25366));
    InMux I__5388 (
            .O(N__25369),
            .I(N__25363));
    LocalMux I__5387 (
            .O(N__25366),
            .I(N__25358));
    LocalMux I__5386 (
            .O(N__25363),
            .I(N__25358));
    Span4Mux_h I__5385 (
            .O(N__25358),
            .I(N__25355));
    Odrv4 I__5384 (
            .O(N__25355),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_1 ));
    InMux I__5383 (
            .O(N__25352),
            .I(N__25349));
    LocalMux I__5382 (
            .O(N__25349),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1 ));
    CEMux I__5381 (
            .O(N__25346),
            .I(N__25343));
    LocalMux I__5380 (
            .O(N__25343),
            .I(N__25340));
    Span4Mux_h I__5379 (
            .O(N__25340),
            .I(N__25336));
    CEMux I__5378 (
            .O(N__25339),
            .I(N__25331));
    Span4Mux_v I__5377 (
            .O(N__25336),
            .I(N__25328));
    CEMux I__5376 (
            .O(N__25335),
            .I(N__25325));
    CEMux I__5375 (
            .O(N__25334),
            .I(N__25322));
    LocalMux I__5374 (
            .O(N__25331),
            .I(N__25319));
    Span4Mux_v I__5373 (
            .O(N__25328),
            .I(N__25314));
    LocalMux I__5372 (
            .O(N__25325),
            .I(N__25314));
    LocalMux I__5371 (
            .O(N__25322),
            .I(N__25311));
    Span4Mux_v I__5370 (
            .O(N__25319),
            .I(N__25308));
    Span4Mux_v I__5369 (
            .O(N__25314),
            .I(N__25305));
    Sp12to4 I__5368 (
            .O(N__25311),
            .I(N__25302));
    Span4Mux_s0_h I__5367 (
            .O(N__25308),
            .I(N__25299));
    IoSpan4Mux I__5366 (
            .O(N__25305),
            .I(N__25296));
    Span12Mux_v I__5365 (
            .O(N__25302),
            .I(N__25291));
    Sp12to4 I__5364 (
            .O(N__25299),
            .I(N__25291));
    Span4Mux_s3_v I__5363 (
            .O(N__25296),
            .I(N__25288));
    Odrv12 I__5362 (
            .O(N__25291),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0 ));
    Odrv4 I__5361 (
            .O(N__25288),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0 ));
    InMux I__5360 (
            .O(N__25283),
            .I(N__25279));
    InMux I__5359 (
            .O(N__25282),
            .I(N__25276));
    LocalMux I__5358 (
            .O(N__25279),
            .I(N__25273));
    LocalMux I__5357 (
            .O(N__25276),
            .I(N__25270));
    Span4Mux_h I__5356 (
            .O(N__25273),
            .I(N__25265));
    Span4Mux_s3_h I__5355 (
            .O(N__25270),
            .I(N__25265));
    Odrv4 I__5354 (
            .O(N__25265),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_4 ));
    CascadeMux I__5353 (
            .O(N__25262),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_4_cascade_ ));
    InMux I__5352 (
            .O(N__25259),
            .I(N__25256));
    LocalMux I__5351 (
            .O(N__25256),
            .I(N__25253));
    Span4Mux_v I__5350 (
            .O(N__25253),
            .I(N__25249));
    InMux I__5349 (
            .O(N__25252),
            .I(N__25246));
    Odrv4 I__5348 (
            .O(N__25249),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4 ));
    LocalMux I__5347 (
            .O(N__25246),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4 ));
    CascadeMux I__5346 (
            .O(N__25241),
            .I(N__25238));
    InMux I__5345 (
            .O(N__25238),
            .I(N__25234));
    CascadeMux I__5344 (
            .O(N__25237),
            .I(N__25231));
    LocalMux I__5343 (
            .O(N__25234),
            .I(N__25228));
    InMux I__5342 (
            .O(N__25231),
            .I(N__25225));
    Odrv12 I__5341 (
            .O(N__25228),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4 ));
    LocalMux I__5340 (
            .O(N__25225),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4 ));
    InMux I__5339 (
            .O(N__25220),
            .I(N__25217));
    LocalMux I__5338 (
            .O(N__25217),
            .I(N__25213));
    InMux I__5337 (
            .O(N__25216),
            .I(N__25210));
    Span4Mux_v I__5336 (
            .O(N__25213),
            .I(N__25205));
    LocalMux I__5335 (
            .O(N__25210),
            .I(N__25205));
    Span4Mux_v I__5334 (
            .O(N__25205),
            .I(N__25202));
    Span4Mux_s1_v I__5333 (
            .O(N__25202),
            .I(N__25199));
    Odrv4 I__5332 (
            .O(N__25199),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_4 ));
    InMux I__5331 (
            .O(N__25196),
            .I(N__25192));
    InMux I__5330 (
            .O(N__25195),
            .I(N__25189));
    LocalMux I__5329 (
            .O(N__25192),
            .I(N__25186));
    LocalMux I__5328 (
            .O(N__25189),
            .I(N__25183));
    Span12Mux_v I__5327 (
            .O(N__25186),
            .I(N__25180));
    Span4Mux_h I__5326 (
            .O(N__25183),
            .I(N__25177));
    Odrv12 I__5325 (
            .O(N__25180),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4 ));
    Odrv4 I__5324 (
            .O(N__25177),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4 ));
    CascadeMux I__5323 (
            .O(N__25172),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_4_cascade_ ));
    InMux I__5322 (
            .O(N__25169),
            .I(N__25166));
    LocalMux I__5321 (
            .O(N__25166),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_4 ));
    CascadeMux I__5320 (
            .O(N__25163),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_4_cascade_ ));
    CascadeMux I__5319 (
            .O(N__25160),
            .I(N__25157));
    InMux I__5318 (
            .O(N__25157),
            .I(N__25154));
    LocalMux I__5317 (
            .O(N__25154),
            .I(N__25151));
    Odrv12 I__5316 (
            .O(N__25151),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_4 ));
    CascadeMux I__5315 (
            .O(N__25148),
            .I(N__25144));
    InMux I__5314 (
            .O(N__25147),
            .I(N__25139));
    InMux I__5313 (
            .O(N__25144),
            .I(N__25139));
    LocalMux I__5312 (
            .O(N__25139),
            .I(N__25136));
    Odrv4 I__5311 (
            .O(N__25136),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_4 ));
    CascadeMux I__5310 (
            .O(N__25133),
            .I(N__25130));
    InMux I__5309 (
            .O(N__25130),
            .I(N__25124));
    InMux I__5308 (
            .O(N__25129),
            .I(N__25124));
    LocalMux I__5307 (
            .O(N__25124),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_4 ));
    CascadeMux I__5306 (
            .O(N__25121),
            .I(N__25118));
    InMux I__5305 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__5304 (
            .O(N__25115),
            .I(N__25112));
    Odrv4 I__5303 (
            .O(N__25112),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_4 ));
    InMux I__5302 (
            .O(N__25109),
            .I(N__25105));
    InMux I__5301 (
            .O(N__25108),
            .I(N__25102));
    LocalMux I__5300 (
            .O(N__25105),
            .I(N__25097));
    LocalMux I__5299 (
            .O(N__25102),
            .I(N__25097));
    Span4Mux_h I__5298 (
            .O(N__25097),
            .I(N__25094));
    Odrv4 I__5297 (
            .O(N__25094),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_4 ));
    CEMux I__5296 (
            .O(N__25091),
            .I(N__25088));
    LocalMux I__5295 (
            .O(N__25088),
            .I(N__25084));
    CEMux I__5294 (
            .O(N__25087),
            .I(N__25081));
    Span4Mux_v I__5293 (
            .O(N__25084),
            .I(N__25078));
    LocalMux I__5292 (
            .O(N__25081),
            .I(N__25075));
    Span4Mux_h I__5291 (
            .O(N__25078),
            .I(N__25072));
    Span4Mux_v I__5290 (
            .O(N__25075),
            .I(N__25069));
    Sp12to4 I__5289 (
            .O(N__25072),
            .I(N__25064));
    Sp12to4 I__5288 (
            .O(N__25069),
            .I(N__25064));
    Odrv12 I__5287 (
            .O(N__25064),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe16 ));
    InMux I__5286 (
            .O(N__25061),
            .I(N__25058));
    LocalMux I__5285 (
            .O(N__25058),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1 ));
    CascadeMux I__5284 (
            .O(N__25055),
            .I(N__25052));
    InMux I__5283 (
            .O(N__25052),
            .I(N__25049));
    LocalMux I__5282 (
            .O(N__25049),
            .I(N__25045));
    InMux I__5281 (
            .O(N__25048),
            .I(N__25042));
    Span4Mux_h I__5280 (
            .O(N__25045),
            .I(N__25039));
    LocalMux I__5279 (
            .O(N__25042),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5 ));
    Odrv4 I__5278 (
            .O(N__25039),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5 ));
    InMux I__5277 (
            .O(N__25034),
            .I(N__25030));
    CascadeMux I__5276 (
            .O(N__25033),
            .I(N__25027));
    LocalMux I__5275 (
            .O(N__25030),
            .I(N__25024));
    InMux I__5274 (
            .O(N__25027),
            .I(N__25021));
    Span4Mux_v I__5273 (
            .O(N__25024),
            .I(N__25018));
    LocalMux I__5272 (
            .O(N__25021),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5 ));
    Odrv4 I__5271 (
            .O(N__25018),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5 ));
    CascadeMux I__5270 (
            .O(N__25013),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_5_cascade_ ));
    InMux I__5269 (
            .O(N__25010),
            .I(N__25007));
    LocalMux I__5268 (
            .O(N__25007),
            .I(N__25004));
    Span4Mux_s3_h I__5267 (
            .O(N__25004),
            .I(N__25001));
    Span4Mux_v I__5266 (
            .O(N__25001),
            .I(N__24998));
    Odrv4 I__5265 (
            .O(N__24998),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_5 ));
    InMux I__5264 (
            .O(N__24995),
            .I(N__24992));
    LocalMux I__5263 (
            .O(N__24992),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_5 ));
    CascadeMux I__5262 (
            .O(N__24989),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_5_cascade_ ));
    InMux I__5261 (
            .O(N__24986),
            .I(N__24983));
    LocalMux I__5260 (
            .O(N__24983),
            .I(N__24980));
    Span4Mux_h I__5259 (
            .O(N__24980),
            .I(N__24977));
    Span4Mux_h I__5258 (
            .O(N__24977),
            .I(N__24974));
    Odrv4 I__5257 (
            .O(N__24974),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_5 ));
    InMux I__5256 (
            .O(N__24971),
            .I(N__24968));
    LocalMux I__5255 (
            .O(N__24968),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_1 ));
    InMux I__5254 (
            .O(N__24965),
            .I(N__24962));
    LocalMux I__5253 (
            .O(N__24962),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_1 ));
    InMux I__5252 (
            .O(N__24959),
            .I(N__24956));
    LocalMux I__5251 (
            .O(N__24956),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_1 ));
    InMux I__5250 (
            .O(N__24953),
            .I(N__24947));
    InMux I__5249 (
            .O(N__24952),
            .I(N__24947));
    LocalMux I__5248 (
            .O(N__24947),
            .I(N__24944));
    Odrv4 I__5247 (
            .O(N__24944),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_4 ));
    CascadeMux I__5246 (
            .O(N__24941),
            .I(N__24937));
    InMux I__5245 (
            .O(N__24940),
            .I(N__24934));
    InMux I__5244 (
            .O(N__24937),
            .I(N__24931));
    LocalMux I__5243 (
            .O(N__24934),
            .I(N__24928));
    LocalMux I__5242 (
            .O(N__24931),
            .I(N__24925));
    Span4Mux_v I__5241 (
            .O(N__24928),
            .I(N__24922));
    Odrv4 I__5240 (
            .O(N__24925),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5 ));
    Odrv4 I__5239 (
            .O(N__24922),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5 ));
    CEMux I__5238 (
            .O(N__24917),
            .I(N__24913));
    CEMux I__5237 (
            .O(N__24916),
            .I(N__24910));
    LocalMux I__5236 (
            .O(N__24913),
            .I(N__24907));
    LocalMux I__5235 (
            .O(N__24910),
            .I(N__24904));
    Span4Mux_s2_v I__5234 (
            .O(N__24907),
            .I(N__24901));
    Span12Mux_s8_h I__5233 (
            .O(N__24904),
            .I(N__24898));
    Span4Mux_h I__5232 (
            .O(N__24901),
            .I(N__24895));
    Odrv12 I__5231 (
            .O(N__24898),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17 ));
    Odrv4 I__5230 (
            .O(N__24895),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17 ));
    CascadeMux I__5229 (
            .O(N__24890),
            .I(N__24887));
    InMux I__5228 (
            .O(N__24887),
            .I(N__24884));
    LocalMux I__5227 (
            .O(N__24884),
            .I(N__24881));
    Span4Mux_v I__5226 (
            .O(N__24881),
            .I(N__24878));
    Span4Mux_s3_h I__5225 (
            .O(N__24878),
            .I(N__24874));
    InMux I__5224 (
            .O(N__24877),
            .I(N__24871));
    Odrv4 I__5223 (
            .O(N__24874),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6 ));
    LocalMux I__5222 (
            .O(N__24871),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6 ));
    InMux I__5221 (
            .O(N__24866),
            .I(N__24863));
    LocalMux I__5220 (
            .O(N__24863),
            .I(N__24859));
    InMux I__5219 (
            .O(N__24862),
            .I(N__24856));
    Span4Mux_v I__5218 (
            .O(N__24859),
            .I(N__24851));
    LocalMux I__5217 (
            .O(N__24856),
            .I(N__24851));
    Span4Mux_v I__5216 (
            .O(N__24851),
            .I(N__24848));
    Odrv4 I__5215 (
            .O(N__24848),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_6 ));
    InMux I__5214 (
            .O(N__24845),
            .I(N__24842));
    LocalMux I__5213 (
            .O(N__24842),
            .I(N__24839));
    Odrv12 I__5212 (
            .O(N__24839),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_6 ));
    CascadeMux I__5211 (
            .O(N__24836),
            .I(N__24833));
    InMux I__5210 (
            .O(N__24833),
            .I(N__24829));
    CascadeMux I__5209 (
            .O(N__24832),
            .I(N__24826));
    LocalMux I__5208 (
            .O(N__24829),
            .I(N__24823));
    InMux I__5207 (
            .O(N__24826),
            .I(N__24820));
    Odrv4 I__5206 (
            .O(N__24823),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0 ));
    LocalMux I__5205 (
            .O(N__24820),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0 ));
    CascadeMux I__5204 (
            .O(N__24815),
            .I(N__24812));
    InMux I__5203 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__5202 (
            .O(N__24809),
            .I(N__24805));
    InMux I__5201 (
            .O(N__24808),
            .I(N__24802));
    Span4Mux_v I__5200 (
            .O(N__24805),
            .I(N__24799));
    LocalMux I__5199 (
            .O(N__24802),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0 ));
    Odrv4 I__5198 (
            .O(N__24799),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0 ));
    CascadeMux I__5197 (
            .O(N__24794),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_0_cascade_ ));
    CascadeMux I__5196 (
            .O(N__24791),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI86UU1_0_cascade_ ));
    InMux I__5195 (
            .O(N__24788),
            .I(N__24785));
    LocalMux I__5194 (
            .O(N__24785),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNI2KHQ1_0 ));
    CascadeMux I__5193 (
            .O(N__24782),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_0_cascade_ ));
    InMux I__5192 (
            .O(N__24779),
            .I(N__24776));
    LocalMux I__5191 (
            .O(N__24776),
            .I(N__24773));
    Span4Mux_v I__5190 (
            .O(N__24773),
            .I(N__24770));
    Span4Mux_h I__5189 (
            .O(N__24770),
            .I(N__24767));
    Odrv4 I__5188 (
            .O(N__24767),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFG9I8_0 ));
    InMux I__5187 (
            .O(N__24764),
            .I(N__24761));
    LocalMux I__5186 (
            .O(N__24761),
            .I(N__24757));
    InMux I__5185 (
            .O(N__24760),
            .I(N__24754));
    Span4Mux_s3_h I__5184 (
            .O(N__24757),
            .I(N__24751));
    LocalMux I__5183 (
            .O(N__24754),
            .I(N__24748));
    Odrv4 I__5182 (
            .O(N__24751),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0 ));
    Odrv12 I__5181 (
            .O(N__24748),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0 ));
    CascadeMux I__5180 (
            .O(N__24743),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_0_cascade_ ));
    InMux I__5179 (
            .O(N__24740),
            .I(N__24737));
    LocalMux I__5178 (
            .O(N__24737),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIKPJ32_0 ));
    InMux I__5177 (
            .O(N__24734),
            .I(N__24731));
    LocalMux I__5176 (
            .O(N__24731),
            .I(N__24728));
    Odrv4 I__5175 (
            .O(N__24728),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_0 ));
    InMux I__5174 (
            .O(N__24725),
            .I(N__24722));
    LocalMux I__5173 (
            .O(N__24722),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI4QLM1_0 ));
    InMux I__5172 (
            .O(N__24719),
            .I(N__24715));
    InMux I__5171 (
            .O(N__24718),
            .I(N__24712));
    LocalMux I__5170 (
            .O(N__24715),
            .I(N__24709));
    LocalMux I__5169 (
            .O(N__24712),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0 ));
    Odrv12 I__5168 (
            .O(N__24709),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0 ));
    CascadeMux I__5167 (
            .O(N__24704),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_0_cascade_ ));
    InMux I__5166 (
            .O(N__24701),
            .I(N__24698));
    LocalMux I__5165 (
            .O(N__24698),
            .I(N__24695));
    Odrv4 I__5164 (
            .O(N__24695),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_0 ));
    CascadeMux I__5163 (
            .O(N__24692),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_0_cascade_ ));
    InMux I__5162 (
            .O(N__24689),
            .I(N__24686));
    LocalMux I__5161 (
            .O(N__24686),
            .I(N__24683));
    Odrv4 I__5160 (
            .O(N__24683),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_0 ));
    InMux I__5159 (
            .O(N__24680),
            .I(N__24677));
    LocalMux I__5158 (
            .O(N__24677),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_0 ));
    InMux I__5157 (
            .O(N__24674),
            .I(N__24671));
    LocalMux I__5156 (
            .O(N__24671),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_0 ));
    InMux I__5155 (
            .O(N__24668),
            .I(N__24662));
    InMux I__5154 (
            .O(N__24667),
            .I(N__24662));
    LocalMux I__5153 (
            .O(N__24662),
            .I(N__24659));
    Odrv12 I__5152 (
            .O(N__24659),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_0 ));
    InMux I__5151 (
            .O(N__24656),
            .I(N__24653));
    LocalMux I__5150 (
            .O(N__24653),
            .I(N__24649));
    InMux I__5149 (
            .O(N__24652),
            .I(N__24646));
    Odrv4 I__5148 (
            .O(N__24649),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0 ));
    LocalMux I__5147 (
            .O(N__24646),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0 ));
    CascadeMux I__5146 (
            .O(N__24641),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_0_cascade_ ));
    InMux I__5145 (
            .O(N__24638),
            .I(N__24635));
    LocalMux I__5144 (
            .O(N__24635),
            .I(N__24632));
    Span4Mux_v I__5143 (
            .O(N__24632),
            .I(N__24628));
    InMux I__5142 (
            .O(N__24631),
            .I(N__24625));
    Odrv4 I__5141 (
            .O(N__24628),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0 ));
    LocalMux I__5140 (
            .O(N__24625),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0 ));
    InMux I__5139 (
            .O(N__24620),
            .I(N__24617));
    LocalMux I__5138 (
            .O(N__24617),
            .I(N__24614));
    Odrv4 I__5137 (
            .O(N__24614),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_6 ));
    InMux I__5136 (
            .O(N__24611),
            .I(N__24608));
    LocalMux I__5135 (
            .O(N__24608),
            .I(N__24605));
    Span4Mux_h I__5134 (
            .O(N__24605),
            .I(N__24602));
    Span4Mux_h I__5133 (
            .O(N__24602),
            .I(N__24599));
    Odrv4 I__5132 (
            .O(N__24599),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_6 ));
    CascadeMux I__5131 (
            .O(N__24596),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_4_cascade_ ));
    CascadeMux I__5130 (
            .O(N__24593),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_4_cascade_ ));
    CascadeMux I__5129 (
            .O(N__24590),
            .I(N__24587));
    InMux I__5128 (
            .O(N__24587),
            .I(N__24584));
    LocalMux I__5127 (
            .O(N__24584),
            .I(N__24581));
    Span4Mux_v I__5126 (
            .O(N__24581),
            .I(N__24578));
    Span4Mux_h I__5125 (
            .O(N__24578),
            .I(N__24575));
    Odrv4 I__5124 (
            .O(N__24575),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_4 ));
    InMux I__5123 (
            .O(N__24572),
            .I(N__24568));
    CascadeMux I__5122 (
            .O(N__24571),
            .I(N__24565));
    LocalMux I__5121 (
            .O(N__24568),
            .I(N__24562));
    InMux I__5120 (
            .O(N__24565),
            .I(N__24559));
    Span4Mux_s3_v I__5119 (
            .O(N__24562),
            .I(N__24554));
    LocalMux I__5118 (
            .O(N__24559),
            .I(N__24554));
    Span4Mux_v I__5117 (
            .O(N__24554),
            .I(N__24551));
    Odrv4 I__5116 (
            .O(N__24551),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_6 ));
    InMux I__5115 (
            .O(N__24548),
            .I(N__24544));
    InMux I__5114 (
            .O(N__24547),
            .I(N__24541));
    LocalMux I__5113 (
            .O(N__24544),
            .I(N__24538));
    LocalMux I__5112 (
            .O(N__24541),
            .I(N__24535));
    Odrv4 I__5111 (
            .O(N__24538),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6 ));
    Odrv12 I__5110 (
            .O(N__24535),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6 ));
    CascadeMux I__5109 (
            .O(N__24530),
            .I(N__24527));
    InMux I__5108 (
            .O(N__24527),
            .I(N__24524));
    LocalMux I__5107 (
            .O(N__24524),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_6 ));
    InMux I__5106 (
            .O(N__24521),
            .I(N__24518));
    LocalMux I__5105 (
            .O(N__24518),
            .I(N__24514));
    InMux I__5104 (
            .O(N__24517),
            .I(N__24511));
    Span4Mux_v I__5103 (
            .O(N__24514),
            .I(N__24508));
    LocalMux I__5102 (
            .O(N__24511),
            .I(N__24505));
    Odrv4 I__5101 (
            .O(N__24508),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4 ));
    Odrv4 I__5100 (
            .O(N__24505),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4 ));
    InMux I__5099 (
            .O(N__24500),
            .I(N__24496));
    InMux I__5098 (
            .O(N__24499),
            .I(N__24493));
    LocalMux I__5097 (
            .O(N__24496),
            .I(N__24490));
    LocalMux I__5096 (
            .O(N__24493),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4 ));
    Odrv4 I__5095 (
            .O(N__24490),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4 ));
    CascadeMux I__5094 (
            .O(N__24485),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_4_cascade_ ));
    InMux I__5093 (
            .O(N__24482),
            .I(N__24479));
    LocalMux I__5092 (
            .O(N__24479),
            .I(N__24475));
    InMux I__5091 (
            .O(N__24478),
            .I(N__24472));
    Odrv4 I__5090 (
            .O(N__24475),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4 ));
    LocalMux I__5089 (
            .O(N__24472),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4 ));
    InMux I__5088 (
            .O(N__24467),
            .I(N__24464));
    LocalMux I__5087 (
            .O(N__24464),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_4 ));
    InMux I__5086 (
            .O(N__24461),
            .I(N__24458));
    LocalMux I__5085 (
            .O(N__24458),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_6 ));
    InMux I__5084 (
            .O(N__24455),
            .I(N__24452));
    LocalMux I__5083 (
            .O(N__24452),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_6 ));
    CascadeMux I__5082 (
            .O(N__24449),
            .I(N__24446));
    InMux I__5081 (
            .O(N__24446),
            .I(N__24440));
    InMux I__5080 (
            .O(N__24445),
            .I(N__24440));
    LocalMux I__5079 (
            .O(N__24440),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_6 ));
    CEMux I__5078 (
            .O(N__24437),
            .I(N__24434));
    LocalMux I__5077 (
            .O(N__24434),
            .I(N__24431));
    Span4Mux_h I__5076 (
            .O(N__24431),
            .I(N__24428));
    Odrv4 I__5075 (
            .O(N__24428),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe28 ));
    InMux I__5074 (
            .O(N__24425),
            .I(N__24421));
    InMux I__5073 (
            .O(N__24424),
            .I(N__24418));
    LocalMux I__5072 (
            .O(N__24421),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5 ));
    LocalMux I__5071 (
            .O(N__24418),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5 ));
    CEMux I__5070 (
            .O(N__24413),
            .I(N__24410));
    LocalMux I__5069 (
            .O(N__24410),
            .I(N__24405));
    CEMux I__5068 (
            .O(N__24409),
            .I(N__24402));
    CEMux I__5067 (
            .O(N__24408),
            .I(N__24399));
    Span4Mux_s3_v I__5066 (
            .O(N__24405),
            .I(N__24394));
    LocalMux I__5065 (
            .O(N__24402),
            .I(N__24394));
    LocalMux I__5064 (
            .O(N__24399),
            .I(N__24391));
    Span4Mux_v I__5063 (
            .O(N__24394),
            .I(N__24388));
    Span4Mux_v I__5062 (
            .O(N__24391),
            .I(N__24385));
    Span4Mux_h I__5061 (
            .O(N__24388),
            .I(N__24382));
    Odrv4 I__5060 (
            .O(N__24385),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30 ));
    Odrv4 I__5059 (
            .O(N__24382),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30 ));
    InMux I__5058 (
            .O(N__24377),
            .I(N__24374));
    LocalMux I__5057 (
            .O(N__24374),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_6 ));
    InMux I__5056 (
            .O(N__24371),
            .I(N__24368));
    LocalMux I__5055 (
            .O(N__24368),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_6 ));
    CascadeMux I__5054 (
            .O(N__24365),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_6_cascade_ ));
    InMux I__5053 (
            .O(N__24362),
            .I(N__24359));
    LocalMux I__5052 (
            .O(N__24359),
            .I(N__24356));
    Odrv4 I__5051 (
            .O(N__24356),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNISIMM1_6 ));
    CascadeMux I__5050 (
            .O(N__24353),
            .I(N__24349));
    InMux I__5049 (
            .O(N__24352),
            .I(N__24344));
    InMux I__5048 (
            .O(N__24349),
            .I(N__24344));
    LocalMux I__5047 (
            .O(N__24344),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_5 ));
    CascadeMux I__5046 (
            .O(N__24341),
            .I(N__24334));
    CascadeMux I__5045 (
            .O(N__24340),
            .I(N__24328));
    CascadeMux I__5044 (
            .O(N__24339),
            .I(N__24324));
    CascadeMux I__5043 (
            .O(N__24338),
            .I(N__24320));
    InMux I__5042 (
            .O(N__24337),
            .I(N__24311));
    InMux I__5041 (
            .O(N__24334),
            .I(N__24301));
    InMux I__5040 (
            .O(N__24333),
            .I(N__24301));
    InMux I__5039 (
            .O(N__24332),
            .I(N__24301));
    InMux I__5038 (
            .O(N__24331),
            .I(N__24294));
    InMux I__5037 (
            .O(N__24328),
            .I(N__24294));
    InMux I__5036 (
            .O(N__24327),
            .I(N__24294));
    InMux I__5035 (
            .O(N__24324),
            .I(N__24279));
    InMux I__5034 (
            .O(N__24323),
            .I(N__24279));
    InMux I__5033 (
            .O(N__24320),
            .I(N__24279));
    InMux I__5032 (
            .O(N__24319),
            .I(N__24279));
    InMux I__5031 (
            .O(N__24318),
            .I(N__24272));
    InMux I__5030 (
            .O(N__24317),
            .I(N__24267));
    InMux I__5029 (
            .O(N__24316),
            .I(N__24267));
    InMux I__5028 (
            .O(N__24315),
            .I(N__24264));
    InMux I__5027 (
            .O(N__24314),
            .I(N__24261));
    LocalMux I__5026 (
            .O(N__24311),
            .I(N__24258));
    InMux I__5025 (
            .O(N__24310),
            .I(N__24255));
    InMux I__5024 (
            .O(N__24309),
            .I(N__24250));
    InMux I__5023 (
            .O(N__24308),
            .I(N__24250));
    LocalMux I__5022 (
            .O(N__24301),
            .I(N__24245));
    LocalMux I__5021 (
            .O(N__24294),
            .I(N__24245));
    InMux I__5020 (
            .O(N__24293),
            .I(N__24240));
    InMux I__5019 (
            .O(N__24292),
            .I(N__24240));
    InMux I__5018 (
            .O(N__24291),
            .I(N__24237));
    InMux I__5017 (
            .O(N__24290),
            .I(N__24230));
    InMux I__5016 (
            .O(N__24289),
            .I(N__24230));
    InMux I__5015 (
            .O(N__24288),
            .I(N__24230));
    LocalMux I__5014 (
            .O(N__24279),
            .I(N__24227));
    InMux I__5013 (
            .O(N__24278),
            .I(N__24218));
    InMux I__5012 (
            .O(N__24277),
            .I(N__24218));
    InMux I__5011 (
            .O(N__24276),
            .I(N__24218));
    InMux I__5010 (
            .O(N__24275),
            .I(N__24218));
    LocalMux I__5009 (
            .O(N__24272),
            .I(N__24215));
    LocalMux I__5008 (
            .O(N__24267),
            .I(N__24212));
    LocalMux I__5007 (
            .O(N__24264),
            .I(N__24203));
    LocalMux I__5006 (
            .O(N__24261),
            .I(N__24203));
    Span4Mux_h I__5005 (
            .O(N__24258),
            .I(N__24203));
    LocalMux I__5004 (
            .O(N__24255),
            .I(N__24203));
    LocalMux I__5003 (
            .O(N__24250),
            .I(N__24194));
    Span4Mux_h I__5002 (
            .O(N__24245),
            .I(N__24194));
    LocalMux I__5001 (
            .O(N__24240),
            .I(N__24194));
    LocalMux I__5000 (
            .O(N__24237),
            .I(N__24194));
    LocalMux I__4999 (
            .O(N__24230),
            .I(N__24187));
    Span4Mux_h I__4998 (
            .O(N__24227),
            .I(N__24187));
    LocalMux I__4997 (
            .O(N__24218),
            .I(N__24187));
    Span4Mux_v I__4996 (
            .O(N__24215),
            .I(N__24178));
    Span4Mux_v I__4995 (
            .O(N__24212),
            .I(N__24178));
    Span4Mux_v I__4994 (
            .O(N__24203),
            .I(N__24178));
    Span4Mux_v I__4993 (
            .O(N__24194),
            .I(N__24178));
    Odrv4 I__4992 (
            .O(N__24187),
            .I(instruction_16));
    Odrv4 I__4991 (
            .O(N__24178),
            .I(instruction_16));
    InMux I__4990 (
            .O(N__24173),
            .I(N__24156));
    InMux I__4989 (
            .O(N__24172),
            .I(N__24156));
    InMux I__4988 (
            .O(N__24171),
            .I(N__24148));
    InMux I__4987 (
            .O(N__24170),
            .I(N__24148));
    CascadeMux I__4986 (
            .O(N__24169),
            .I(N__24144));
    InMux I__4985 (
            .O(N__24168),
            .I(N__24139));
    InMux I__4984 (
            .O(N__24167),
            .I(N__24139));
    InMux I__4983 (
            .O(N__24166),
            .I(N__24136));
    InMux I__4982 (
            .O(N__24165),
            .I(N__24127));
    InMux I__4981 (
            .O(N__24164),
            .I(N__24127));
    InMux I__4980 (
            .O(N__24163),
            .I(N__24127));
    InMux I__4979 (
            .O(N__24162),
            .I(N__24127));
    InMux I__4978 (
            .O(N__24161),
            .I(N__24123));
    LocalMux I__4977 (
            .O(N__24156),
            .I(N__24120));
    InMux I__4976 (
            .O(N__24155),
            .I(N__24113));
    InMux I__4975 (
            .O(N__24154),
            .I(N__24113));
    InMux I__4974 (
            .O(N__24153),
            .I(N__24113));
    LocalMux I__4973 (
            .O(N__24148),
            .I(N__24108));
    InMux I__4972 (
            .O(N__24147),
            .I(N__24105));
    InMux I__4971 (
            .O(N__24144),
            .I(N__24102));
    LocalMux I__4970 (
            .O(N__24139),
            .I(N__24091));
    LocalMux I__4969 (
            .O(N__24136),
            .I(N__24086));
    LocalMux I__4968 (
            .O(N__24127),
            .I(N__24086));
    InMux I__4967 (
            .O(N__24126),
            .I(N__24083));
    LocalMux I__4966 (
            .O(N__24123),
            .I(N__24076));
    Span4Mux_s3_v I__4965 (
            .O(N__24120),
            .I(N__24076));
    LocalMux I__4964 (
            .O(N__24113),
            .I(N__24076));
    InMux I__4963 (
            .O(N__24112),
            .I(N__24073));
    InMux I__4962 (
            .O(N__24111),
            .I(N__24070));
    Span4Mux_v I__4961 (
            .O(N__24108),
            .I(N__24063));
    LocalMux I__4960 (
            .O(N__24105),
            .I(N__24063));
    LocalMux I__4959 (
            .O(N__24102),
            .I(N__24063));
    InMux I__4958 (
            .O(N__24101),
            .I(N__24054));
    InMux I__4957 (
            .O(N__24100),
            .I(N__24054));
    InMux I__4956 (
            .O(N__24099),
            .I(N__24054));
    InMux I__4955 (
            .O(N__24098),
            .I(N__24054));
    InMux I__4954 (
            .O(N__24097),
            .I(N__24045));
    InMux I__4953 (
            .O(N__24096),
            .I(N__24045));
    InMux I__4952 (
            .O(N__24095),
            .I(N__24045));
    InMux I__4951 (
            .O(N__24094),
            .I(N__24045));
    Span4Mux_s3_v I__4950 (
            .O(N__24091),
            .I(N__24036));
    Span4Mux_v I__4949 (
            .O(N__24086),
            .I(N__24036));
    LocalMux I__4948 (
            .O(N__24083),
            .I(N__24036));
    Span4Mux_h I__4947 (
            .O(N__24076),
            .I(N__24036));
    LocalMux I__4946 (
            .O(N__24073),
            .I(N__24025));
    LocalMux I__4945 (
            .O(N__24070),
            .I(N__24025));
    Sp12to4 I__4944 (
            .O(N__24063),
            .I(N__24025));
    LocalMux I__4943 (
            .O(N__24054),
            .I(N__24025));
    LocalMux I__4942 (
            .O(N__24045),
            .I(N__24025));
    Span4Mux_h I__4941 (
            .O(N__24036),
            .I(N__24022));
    Span12Mux_s9_h I__4940 (
            .O(N__24025),
            .I(N__24019));
    Odrv4 I__4939 (
            .O(N__24022),
            .I(instruction_15));
    Odrv12 I__4938 (
            .O(N__24019),
            .I(instruction_15));
    CascadeMux I__4937 (
            .O(N__24014),
            .I(N__24009));
    InMux I__4936 (
            .O(N__24013),
            .I(N__24006));
    InMux I__4935 (
            .O(N__24012),
            .I(N__24003));
    InMux I__4934 (
            .O(N__24009),
            .I(N__24000));
    LocalMux I__4933 (
            .O(N__24006),
            .I(N__23994));
    LocalMux I__4932 (
            .O(N__24003),
            .I(N__23994));
    LocalMux I__4931 (
            .O(N__24000),
            .I(N__23991));
    InMux I__4930 (
            .O(N__23999),
            .I(N__23982));
    Span4Mux_v I__4929 (
            .O(N__23994),
            .I(N__23977));
    Span4Mux_v I__4928 (
            .O(N__23991),
            .I(N__23977));
    InMux I__4927 (
            .O(N__23990),
            .I(N__23971));
    InMux I__4926 (
            .O(N__23989),
            .I(N__23971));
    InMux I__4925 (
            .O(N__23988),
            .I(N__23968));
    InMux I__4924 (
            .O(N__23987),
            .I(N__23965));
    InMux I__4923 (
            .O(N__23986),
            .I(N__23962));
    InMux I__4922 (
            .O(N__23985),
            .I(N__23959));
    LocalMux I__4921 (
            .O(N__23982),
            .I(N__23956));
    IoSpan4Mux I__4920 (
            .O(N__23977),
            .I(N__23953));
    InMux I__4919 (
            .O(N__23976),
            .I(N__23950));
    LocalMux I__4918 (
            .O(N__23971),
            .I(N__23947));
    LocalMux I__4917 (
            .O(N__23968),
            .I(N__23944));
    LocalMux I__4916 (
            .O(N__23965),
            .I(N__23941));
    LocalMux I__4915 (
            .O(N__23962),
            .I(N__23938));
    LocalMux I__4914 (
            .O(N__23959),
            .I(N__23935));
    Span4Mux_v I__4913 (
            .O(N__23956),
            .I(N__23932));
    Span4Mux_s3_h I__4912 (
            .O(N__23953),
            .I(N__23927));
    LocalMux I__4911 (
            .O(N__23950),
            .I(N__23927));
    Span4Mux_v I__4910 (
            .O(N__23947),
            .I(N__23922));
    Span4Mux_h I__4909 (
            .O(N__23944),
            .I(N__23922));
    Span4Mux_h I__4908 (
            .O(N__23941),
            .I(N__23919));
    Span12Mux_s7_h I__4907 (
            .O(N__23938),
            .I(N__23916));
    Span4Mux_h I__4906 (
            .O(N__23935),
            .I(N__23913));
    Span4Mux_h I__4905 (
            .O(N__23932),
            .I(N__23908));
    Span4Mux_h I__4904 (
            .O(N__23927),
            .I(N__23908));
    Span4Mux_v I__4903 (
            .O(N__23922),
            .I(N__23905));
    Odrv4 I__4902 (
            .O(N__23919),
            .I(\processor_zipi8.un28_carry_flag_value_1 ));
    Odrv12 I__4901 (
            .O(N__23916),
            .I(\processor_zipi8.un28_carry_flag_value_1 ));
    Odrv4 I__4900 (
            .O(N__23913),
            .I(\processor_zipi8.un28_carry_flag_value_1 ));
    Odrv4 I__4899 (
            .O(N__23908),
            .I(\processor_zipi8.un28_carry_flag_value_1 ));
    Odrv4 I__4898 (
            .O(N__23905),
            .I(\processor_zipi8.un28_carry_flag_value_1 ));
    InMux I__4897 (
            .O(N__23894),
            .I(N__23891));
    LocalMux I__4896 (
            .O(N__23891),
            .I(N__23887));
    InMux I__4895 (
            .O(N__23890),
            .I(N__23884));
    Span4Mux_h I__4894 (
            .O(N__23887),
            .I(N__23879));
    LocalMux I__4893 (
            .O(N__23884),
            .I(N__23879));
    Span4Mux_v I__4892 (
            .O(N__23879),
            .I(N__23876));
    Odrv4 I__4891 (
            .O(N__23876),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_5 ));
    InMux I__4890 (
            .O(N__23873),
            .I(N__23869));
    InMux I__4889 (
            .O(N__23872),
            .I(N__23866));
    LocalMux I__4888 (
            .O(N__23869),
            .I(N__23863));
    LocalMux I__4887 (
            .O(N__23866),
            .I(N__23860));
    Span4Mux_h I__4886 (
            .O(N__23863),
            .I(N__23857));
    Span4Mux_h I__4885 (
            .O(N__23860),
            .I(N__23854));
    Span4Mux_v I__4884 (
            .O(N__23857),
            .I(N__23851));
    Odrv4 I__4883 (
            .O(N__23854),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7 ));
    Odrv4 I__4882 (
            .O(N__23851),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7 ));
    InMux I__4881 (
            .O(N__23846),
            .I(N__23843));
    LocalMux I__4880 (
            .O(N__23843),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_6 ));
    CascadeMux I__4879 (
            .O(N__23840),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_6_cascade_ ));
    InMux I__4878 (
            .O(N__23837),
            .I(N__23834));
    LocalMux I__4877 (
            .O(N__23834),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_6 ));
    CascadeMux I__4876 (
            .O(N__23831),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_6_cascade_ ));
    InMux I__4875 (
            .O(N__23828),
            .I(N__23825));
    LocalMux I__4874 (
            .O(N__23825),
            .I(N__23822));
    Span4Mux_h I__4873 (
            .O(N__23822),
            .I(N__23819));
    Span4Mux_h I__4872 (
            .O(N__23819),
            .I(N__23816));
    Odrv4 I__4871 (
            .O(N__23816),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_6 ));
    CascadeMux I__4870 (
            .O(N__23813),
            .I(N__23810));
    InMux I__4869 (
            .O(N__23810),
            .I(N__23806));
    InMux I__4868 (
            .O(N__23809),
            .I(N__23803));
    LocalMux I__4867 (
            .O(N__23806),
            .I(N__23798));
    LocalMux I__4866 (
            .O(N__23803),
            .I(N__23798));
    Span4Mux_h I__4865 (
            .O(N__23798),
            .I(N__23795));
    Span4Mux_v I__4864 (
            .O(N__23795),
            .I(N__23792));
    Span4Mux_v I__4863 (
            .O(N__23792),
            .I(N__23789));
    Odrv4 I__4862 (
            .O(N__23789),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_6 ));
    CascadeMux I__4861 (
            .O(N__23786),
            .I(N__23783));
    InMux I__4860 (
            .O(N__23783),
            .I(N__23777));
    InMux I__4859 (
            .O(N__23782),
            .I(N__23777));
    LocalMux I__4858 (
            .O(N__23777),
            .I(N__23774));
    Span4Mux_h I__4857 (
            .O(N__23774),
            .I(N__23771));
    Sp12to4 I__4856 (
            .O(N__23771),
            .I(N__23768));
    Span12Mux_v I__4855 (
            .O(N__23768),
            .I(N__23765));
    Odrv12 I__4854 (
            .O(N__23765),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_7 ));
    CEMux I__4853 (
            .O(N__23762),
            .I(N__23759));
    LocalMux I__4852 (
            .O(N__23759),
            .I(N__23756));
    Span4Mux_h I__4851 (
            .O(N__23756),
            .I(N__23753));
    Span4Mux_v I__4850 (
            .O(N__23753),
            .I(N__23750));
    Odrv4 I__4849 (
            .O(N__23750),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe1 ));
    InMux I__4848 (
            .O(N__23747),
            .I(N__23744));
    LocalMux I__4847 (
            .O(N__23744),
            .I(N__23740));
    InMux I__4846 (
            .O(N__23743),
            .I(N__23737));
    Odrv4 I__4845 (
            .O(N__23740),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5 ));
    LocalMux I__4844 (
            .O(N__23737),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5 ));
    CascadeMux I__4843 (
            .O(N__23732),
            .I(N__23729));
    InMux I__4842 (
            .O(N__23729),
            .I(N__23726));
    LocalMux I__4841 (
            .O(N__23726),
            .I(N__23723));
    Span4Mux_s2_v I__4840 (
            .O(N__23723),
            .I(N__23719));
    InMux I__4839 (
            .O(N__23722),
            .I(N__23716));
    Odrv4 I__4838 (
            .O(N__23719),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5 ));
    LocalMux I__4837 (
            .O(N__23716),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5 ));
    InMux I__4836 (
            .O(N__23711),
            .I(N__23708));
    LocalMux I__4835 (
            .O(N__23708),
            .I(N__23705));
    Span4Mux_h I__4834 (
            .O(N__23705),
            .I(N__23701));
    InMux I__4833 (
            .O(N__23704),
            .I(N__23698));
    Odrv4 I__4832 (
            .O(N__23701),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5 ));
    LocalMux I__4831 (
            .O(N__23698),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5 ));
    CascadeMux I__4830 (
            .O(N__23693),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_5_cascade_ ));
    InMux I__4829 (
            .O(N__23690),
            .I(N__23687));
    LocalMux I__4828 (
            .O(N__23687),
            .I(N__23683));
    InMux I__4827 (
            .O(N__23686),
            .I(N__23680));
    Odrv4 I__4826 (
            .O(N__23683),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5 ));
    LocalMux I__4825 (
            .O(N__23680),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5 ));
    CascadeMux I__4824 (
            .O(N__23675),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_5_cascade_ ));
    InMux I__4823 (
            .O(N__23672),
            .I(N__23669));
    LocalMux I__4822 (
            .O(N__23669),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_123 ));
    CascadeMux I__4821 (
            .O(N__23666),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_99_cascade_ ));
    InMux I__4820 (
            .O(N__23663),
            .I(N__23660));
    LocalMux I__4819 (
            .O(N__23660),
            .I(N__23657));
    Span4Mux_s3_h I__4818 (
            .O(N__23657),
            .I(N__23654));
    Span4Mux_h I__4817 (
            .O(N__23654),
            .I(N__23651));
    Odrv4 I__4816 (
            .O(N__23651),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_5 ));
    InMux I__4815 (
            .O(N__23648),
            .I(N__23645));
    LocalMux I__4814 (
            .O(N__23645),
            .I(N__23642));
    Span4Mux_v I__4813 (
            .O(N__23642),
            .I(N__23639));
    Span4Mux_h I__4812 (
            .O(N__23639),
            .I(N__23636));
    Odrv4 I__4811 (
            .O(N__23636),
            .I(\processor_zipi8.stack_memory_3 ));
    InMux I__4810 (
            .O(N__23633),
            .I(N__23630));
    LocalMux I__4809 (
            .O(N__23630),
            .I(N__23627));
    Span4Mux_h I__4808 (
            .O(N__23627),
            .I(N__23624));
    Odrv4 I__4807 (
            .O(N__23624),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_3 ));
    CascadeMux I__4806 (
            .O(N__23621),
            .I(N__23618));
    InMux I__4805 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__4804 (
            .O(N__23615),
            .I(N__23612));
    Span4Mux_v I__4803 (
            .O(N__23612),
            .I(N__23608));
    InMux I__4802 (
            .O(N__23611),
            .I(N__23605));
    Odrv4 I__4801 (
            .O(N__23608),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3 ));
    LocalMux I__4800 (
            .O(N__23605),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3 ));
    InMux I__4799 (
            .O(N__23600),
            .I(N__23597));
    LocalMux I__4798 (
            .O(N__23597),
            .I(N__23593));
    CascadeMux I__4797 (
            .O(N__23596),
            .I(N__23590));
    Span4Mux_s3_v I__4796 (
            .O(N__23593),
            .I(N__23587));
    InMux I__4795 (
            .O(N__23590),
            .I(N__23584));
    Odrv4 I__4794 (
            .O(N__23587),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3 ));
    LocalMux I__4793 (
            .O(N__23584),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3 ));
    InMux I__4792 (
            .O(N__23579),
            .I(N__23576));
    LocalMux I__4791 (
            .O(N__23576),
            .I(N__23573));
    Odrv4 I__4790 (
            .O(N__23573),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_3 ));
    CEMux I__4789 (
            .O(N__23570),
            .I(N__23567));
    LocalMux I__4788 (
            .O(N__23567),
            .I(N__23564));
    Span4Mux_h I__4787 (
            .O(N__23564),
            .I(N__23560));
    CEMux I__4786 (
            .O(N__23563),
            .I(N__23557));
    Span4Mux_s1_h I__4785 (
            .O(N__23560),
            .I(N__23554));
    LocalMux I__4784 (
            .O(N__23557),
            .I(N__23551));
    Sp12to4 I__4783 (
            .O(N__23554),
            .I(N__23548));
    Span4Mux_h I__4782 (
            .O(N__23551),
            .I(N__23545));
    Span12Mux_v I__4781 (
            .O(N__23548),
            .I(N__23542));
    Sp12to4 I__4780 (
            .O(N__23545),
            .I(N__23539));
    Odrv12 I__4779 (
            .O(N__23542),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4 ));
    Odrv12 I__4778 (
            .O(N__23539),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4 ));
    InMux I__4777 (
            .O(N__23534),
            .I(N__23530));
    InMux I__4776 (
            .O(N__23533),
            .I(N__23527));
    LocalMux I__4775 (
            .O(N__23530),
            .I(N__23524));
    LocalMux I__4774 (
            .O(N__23527),
            .I(N__23521));
    Span4Mux_v I__4773 (
            .O(N__23524),
            .I(N__23518));
    Span4Mux_v I__4772 (
            .O(N__23521),
            .I(N__23515));
    Odrv4 I__4771 (
            .O(N__23518),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0 ));
    Odrv4 I__4770 (
            .O(N__23515),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0 ));
    CascadeMux I__4769 (
            .O(N__23510),
            .I(N__23506));
    CascadeMux I__4768 (
            .O(N__23509),
            .I(N__23503));
    InMux I__4767 (
            .O(N__23506),
            .I(N__23500));
    InMux I__4766 (
            .O(N__23503),
            .I(N__23497));
    LocalMux I__4765 (
            .O(N__23500),
            .I(N__23494));
    LocalMux I__4764 (
            .O(N__23497),
            .I(N__23491));
    Odrv4 I__4763 (
            .O(N__23494),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1 ));
    Odrv12 I__4762 (
            .O(N__23491),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1 ));
    CascadeMux I__4761 (
            .O(N__23486),
            .I(N__23482));
    InMux I__4760 (
            .O(N__23485),
            .I(N__23479));
    InMux I__4759 (
            .O(N__23482),
            .I(N__23476));
    LocalMux I__4758 (
            .O(N__23479),
            .I(N__23473));
    LocalMux I__4757 (
            .O(N__23476),
            .I(N__23470));
    Span4Mux_h I__4756 (
            .O(N__23473),
            .I(N__23467));
    Odrv4 I__4755 (
            .O(N__23470),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3 ));
    Odrv4 I__4754 (
            .O(N__23467),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3 ));
    CascadeMux I__4753 (
            .O(N__23462),
            .I(N__23458));
    InMux I__4752 (
            .O(N__23461),
            .I(N__23455));
    InMux I__4751 (
            .O(N__23458),
            .I(N__23452));
    LocalMux I__4750 (
            .O(N__23455),
            .I(N__23447));
    LocalMux I__4749 (
            .O(N__23452),
            .I(N__23447));
    Sp12to4 I__4748 (
            .O(N__23447),
            .I(N__23444));
    Span12Mux_s11_v I__4747 (
            .O(N__23444),
            .I(N__23441));
    Odrv12 I__4746 (
            .O(N__23441),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_6 ));
    CEMux I__4745 (
            .O(N__23438),
            .I(N__23434));
    CEMux I__4744 (
            .O(N__23437),
            .I(N__23431));
    LocalMux I__4743 (
            .O(N__23434),
            .I(N__23428));
    LocalMux I__4742 (
            .O(N__23431),
            .I(N__23425));
    Span4Mux_v I__4741 (
            .O(N__23428),
            .I(N__23422));
    Span4Mux_s0_v I__4740 (
            .O(N__23425),
            .I(N__23419));
    Span4Mux_v I__4739 (
            .O(N__23422),
            .I(N__23416));
    Odrv4 I__4738 (
            .O(N__23419),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5 ));
    Odrv4 I__4737 (
            .O(N__23416),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5 ));
    InMux I__4736 (
            .O(N__23411),
            .I(N__23408));
    LocalMux I__4735 (
            .O(N__23408),
            .I(N__23404));
    InMux I__4734 (
            .O(N__23407),
            .I(N__23401));
    Span4Mux_h I__4733 (
            .O(N__23404),
            .I(N__23398));
    LocalMux I__4732 (
            .O(N__23401),
            .I(N__23395));
    Span4Mux_v I__4731 (
            .O(N__23398),
            .I(N__23390));
    Span4Mux_h I__4730 (
            .O(N__23395),
            .I(N__23390));
    Odrv4 I__4729 (
            .O(N__23390),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_0 ));
    InMux I__4728 (
            .O(N__23387),
            .I(N__23383));
    InMux I__4727 (
            .O(N__23386),
            .I(N__23380));
    LocalMux I__4726 (
            .O(N__23383),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2 ));
    LocalMux I__4725 (
            .O(N__23380),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2 ));
    InMux I__4724 (
            .O(N__23375),
            .I(N__23372));
    LocalMux I__4723 (
            .O(N__23372),
            .I(N__23368));
    InMux I__4722 (
            .O(N__23371),
            .I(N__23365));
    Odrv4 I__4721 (
            .O(N__23368),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2 ));
    LocalMux I__4720 (
            .O(N__23365),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2 ));
    CascadeMux I__4719 (
            .O(N__23360),
            .I(N__23356));
    InMux I__4718 (
            .O(N__23359),
            .I(N__23351));
    InMux I__4717 (
            .O(N__23356),
            .I(N__23351));
    LocalMux I__4716 (
            .O(N__23351),
            .I(N__23348));
    Span4Mux_v I__4715 (
            .O(N__23348),
            .I(N__23345));
    Sp12to4 I__4714 (
            .O(N__23345),
            .I(N__23342));
    Odrv12 I__4713 (
            .O(N__23342),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_4 ));
    InMux I__4712 (
            .O(N__23339),
            .I(N__23335));
    InMux I__4711 (
            .O(N__23338),
            .I(N__23332));
    LocalMux I__4710 (
            .O(N__23335),
            .I(N__23329));
    LocalMux I__4709 (
            .O(N__23332),
            .I(N__23326));
    Span4Mux_v I__4708 (
            .O(N__23329),
            .I(N__23323));
    Span12Mux_s10_v I__4707 (
            .O(N__23326),
            .I(N__23320));
    Odrv4 I__4706 (
            .O(N__23323),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5 ));
    Odrv12 I__4705 (
            .O(N__23320),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5 ));
    InMux I__4704 (
            .O(N__23315),
            .I(N__23312));
    LocalMux I__4703 (
            .O(N__23312),
            .I(N__23308));
    InMux I__4702 (
            .O(N__23311),
            .I(N__23305));
    Span4Mux_v I__4701 (
            .O(N__23308),
            .I(N__23302));
    LocalMux I__4700 (
            .O(N__23305),
            .I(N__23299));
    Span4Mux_v I__4699 (
            .O(N__23302),
            .I(N__23294));
    Span4Mux_v I__4698 (
            .O(N__23299),
            .I(N__23294));
    Odrv4 I__4697 (
            .O(N__23294),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_7 ));
    CEMux I__4696 (
            .O(N__23291),
            .I(N__23288));
    LocalMux I__4695 (
            .O(N__23288),
            .I(N__23285));
    Span4Mux_v I__4694 (
            .O(N__23285),
            .I(N__23282));
    Span4Mux_h I__4693 (
            .O(N__23282),
            .I(N__23279));
    Odrv4 I__4692 (
            .O(N__23279),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe23 ));
    InMux I__4691 (
            .O(N__23276),
            .I(N__23272));
    CascadeMux I__4690 (
            .O(N__23275),
            .I(N__23269));
    LocalMux I__4689 (
            .O(N__23272),
            .I(N__23266));
    InMux I__4688 (
            .O(N__23269),
            .I(N__23263));
    Span4Mux_v I__4687 (
            .O(N__23266),
            .I(N__23258));
    LocalMux I__4686 (
            .O(N__23263),
            .I(N__23258));
    Odrv4 I__4685 (
            .O(N__23258),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_0 ));
    InMux I__4684 (
            .O(N__23255),
            .I(N__23252));
    LocalMux I__4683 (
            .O(N__23252),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_1_0 ));
    InMux I__4682 (
            .O(N__23249),
            .I(N__23245));
    InMux I__4681 (
            .O(N__23248),
            .I(N__23242));
    LocalMux I__4680 (
            .O(N__23245),
            .I(N__23237));
    LocalMux I__4679 (
            .O(N__23242),
            .I(N__23237));
    Span4Mux_v I__4678 (
            .O(N__23237),
            .I(N__23234));
    Odrv4 I__4677 (
            .O(N__23234),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_1 ));
    CascadeMux I__4676 (
            .O(N__23231),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_1_cascade_ ));
    CascadeMux I__4675 (
            .O(N__23228),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_cascade_ ));
    InMux I__4674 (
            .O(N__23225),
            .I(N__23222));
    LocalMux I__4673 (
            .O(N__23222),
            .I(N__23219));
    Odrv4 I__4672 (
            .O(N__23219),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1 ));
    CascadeMux I__4671 (
            .O(N__23216),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_cascade_ ));
    InMux I__4670 (
            .O(N__23213),
            .I(N__23210));
    LocalMux I__4669 (
            .O(N__23210),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1 ));
    CascadeMux I__4668 (
            .O(N__23207),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_cascade_ ));
    InMux I__4667 (
            .O(N__23204),
            .I(N__23201));
    LocalMux I__4666 (
            .O(N__23201),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_1 ));
    InMux I__4665 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__4664 (
            .O(N__23195),
            .I(N__23192));
    Span4Mux_v I__4663 (
            .O(N__23192),
            .I(N__23188));
    InMux I__4662 (
            .O(N__23191),
            .I(N__23185));
    Odrv4 I__4661 (
            .O(N__23188),
            .I(\processor_zipi8.sy_1 ));
    LocalMux I__4660 (
            .O(N__23185),
            .I(\processor_zipi8.sy_1 ));
    CascadeMux I__4659 (
            .O(N__23180),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_4_cascade_ ));
    InMux I__4658 (
            .O(N__23177),
            .I(N__23174));
    LocalMux I__4657 (
            .O(N__23174),
            .I(N__23171));
    Span4Mux_v I__4656 (
            .O(N__23171),
            .I(N__23168));
    Odrv4 I__4655 (
            .O(N__23168),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNICSGN1_4 ));
    CascadeMux I__4654 (
            .O(N__23165),
            .I(N__23160));
    CascadeMux I__4653 (
            .O(N__23164),
            .I(N__23155));
    CascadeMux I__4652 (
            .O(N__23163),
            .I(N__23150));
    InMux I__4651 (
            .O(N__23160),
            .I(N__23147));
    InMux I__4650 (
            .O(N__23159),
            .I(N__23133));
    InMux I__4649 (
            .O(N__23158),
            .I(N__23133));
    InMux I__4648 (
            .O(N__23155),
            .I(N__23133));
    InMux I__4647 (
            .O(N__23154),
            .I(N__23133));
    InMux I__4646 (
            .O(N__23153),
            .I(N__23133));
    InMux I__4645 (
            .O(N__23150),
            .I(N__23133));
    LocalMux I__4644 (
            .O(N__23147),
            .I(N__23130));
    InMux I__4643 (
            .O(N__23146),
            .I(N__23127));
    LocalMux I__4642 (
            .O(N__23133),
            .I(N__23124));
    Span4Mux_h I__4641 (
            .O(N__23130),
            .I(N__23119));
    LocalMux I__4640 (
            .O(N__23127),
            .I(N__23119));
    Span4Mux_v I__4639 (
            .O(N__23124),
            .I(N__23116));
    Span4Mux_v I__4638 (
            .O(N__23119),
            .I(N__23113));
    Odrv4 I__4637 (
            .O(N__23116),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210 ));
    Odrv4 I__4636 (
            .O(N__23113),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210 ));
    CascadeMux I__4635 (
            .O(N__23108),
            .I(N__23100));
    CascadeMux I__4634 (
            .O(N__23107),
            .I(N__23096));
    CascadeMux I__4633 (
            .O(N__23106),
            .I(N__23093));
    CascadeMux I__4632 (
            .O(N__23105),
            .I(N__23089));
    InMux I__4631 (
            .O(N__23104),
            .I(N__23078));
    InMux I__4630 (
            .O(N__23103),
            .I(N__23078));
    InMux I__4629 (
            .O(N__23100),
            .I(N__23078));
    InMux I__4628 (
            .O(N__23099),
            .I(N__23078));
    InMux I__4627 (
            .O(N__23096),
            .I(N__23078));
    InMux I__4626 (
            .O(N__23093),
            .I(N__23071));
    InMux I__4625 (
            .O(N__23092),
            .I(N__23071));
    InMux I__4624 (
            .O(N__23089),
            .I(N__23071));
    LocalMux I__4623 (
            .O(N__23078),
            .I(N__23066));
    LocalMux I__4622 (
            .O(N__23071),
            .I(N__23066));
    Span4Mux_h I__4621 (
            .O(N__23066),
            .I(N__23063));
    Span4Mux_v I__4620 (
            .O(N__23063),
            .I(N__23060));
    Odrv4 I__4619 (
            .O(N__23060),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1211 ));
    CascadeMux I__4618 (
            .O(N__23057),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_0_cascade_ ));
    CascadeMux I__4617 (
            .O(N__23054),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_1_0_cascade_ ));
    InMux I__4616 (
            .O(N__23051),
            .I(N__23048));
    LocalMux I__4615 (
            .O(N__23048),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_0 ));
    CascadeMux I__4614 (
            .O(N__23045),
            .I(N__23042));
    InMux I__4613 (
            .O(N__23042),
            .I(N__23039));
    LocalMux I__4612 (
            .O(N__23039),
            .I(N__23036));
    Span4Mux_h I__4611 (
            .O(N__23036),
            .I(N__23033));
    Span4Mux_v I__4610 (
            .O(N__23033),
            .I(N__23030));
    Odrv4 I__4609 (
            .O(N__23030),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_0 ));
    InMux I__4608 (
            .O(N__23027),
            .I(N__23024));
    LocalMux I__4607 (
            .O(N__23024),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_0 ));
    CascadeMux I__4606 (
            .O(N__23021),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_0_cascade_ ));
    InMux I__4605 (
            .O(N__23018),
            .I(N__23015));
    LocalMux I__4604 (
            .O(N__23015),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_0 ));
    CascadeMux I__4603 (
            .O(N__23012),
            .I(N__23009));
    InMux I__4602 (
            .O(N__23009),
            .I(N__23006));
    LocalMux I__4601 (
            .O(N__23006),
            .I(N__23002));
    InMux I__4600 (
            .O(N__23005),
            .I(N__22999));
    Span4Mux_v I__4599 (
            .O(N__23002),
            .I(N__22996));
    LocalMux I__4598 (
            .O(N__22999),
            .I(N__22993));
    Span4Mux_s1_h I__4597 (
            .O(N__22996),
            .I(N__22990));
    Span4Mux_h I__4596 (
            .O(N__22993),
            .I(N__22987));
    Span4Mux_h I__4595 (
            .O(N__22990),
            .I(N__22984));
    Odrv4 I__4594 (
            .O(N__22987),
            .I(\processor_zipi8.sy_0 ));
    Odrv4 I__4593 (
            .O(N__22984),
            .I(\processor_zipi8.sy_0 ));
    InMux I__4592 (
            .O(N__22979),
            .I(N__22975));
    InMux I__4591 (
            .O(N__22978),
            .I(N__22972));
    LocalMux I__4590 (
            .O(N__22975),
            .I(N__22969));
    LocalMux I__4589 (
            .O(N__22972),
            .I(N__22966));
    Span4Mux_v I__4588 (
            .O(N__22969),
            .I(N__22963));
    Span4Mux_v I__4587 (
            .O(N__22966),
            .I(N__22960));
    Span4Mux_v I__4586 (
            .O(N__22963),
            .I(N__22957));
    Span4Mux_v I__4585 (
            .O(N__22960),
            .I(N__22954));
    Odrv4 I__4584 (
            .O(N__22957),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4 ));
    Odrv4 I__4583 (
            .O(N__22954),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4 ));
    InMux I__4582 (
            .O(N__22949),
            .I(N__22945));
    InMux I__4581 (
            .O(N__22948),
            .I(N__22942));
    LocalMux I__4580 (
            .O(N__22945),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5 ));
    LocalMux I__4579 (
            .O(N__22942),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5 ));
    CEMux I__4578 (
            .O(N__22937),
            .I(N__22934));
    LocalMux I__4577 (
            .O(N__22934),
            .I(N__22931));
    Span4Mux_v I__4576 (
            .O(N__22931),
            .I(N__22927));
    CEMux I__4575 (
            .O(N__22930),
            .I(N__22924));
    Sp12to4 I__4574 (
            .O(N__22927),
            .I(N__22921));
    LocalMux I__4573 (
            .O(N__22924),
            .I(N__22918));
    Odrv12 I__4572 (
            .O(N__22921),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19 ));
    Odrv4 I__4571 (
            .O(N__22918),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19 ));
    InMux I__4570 (
            .O(N__22913),
            .I(N__22910));
    LocalMux I__4569 (
            .O(N__22910),
            .I(N__22906));
    InMux I__4568 (
            .O(N__22909),
            .I(N__22903));
    Odrv12 I__4567 (
            .O(N__22906),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6 ));
    LocalMux I__4566 (
            .O(N__22903),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6 ));
    InMux I__4565 (
            .O(N__22898),
            .I(N__22894));
    InMux I__4564 (
            .O(N__22897),
            .I(N__22891));
    LocalMux I__4563 (
            .O(N__22894),
            .I(N__22888));
    LocalMux I__4562 (
            .O(N__22891),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6 ));
    Odrv12 I__4561 (
            .O(N__22888),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6 ));
    CascadeMux I__4560 (
            .O(N__22883),
            .I(N__22880));
    InMux I__4559 (
            .O(N__22880),
            .I(N__22877));
    LocalMux I__4558 (
            .O(N__22877),
            .I(N__22874));
    Span12Mux_s3_h I__4557 (
            .O(N__22874),
            .I(N__22871));
    Odrv12 I__4556 (
            .O(N__22871),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIUGIQ1_7 ));
    InMux I__4555 (
            .O(N__22868),
            .I(N__22865));
    LocalMux I__4554 (
            .O(N__22865),
            .I(N__22862));
    Span4Mux_h I__4553 (
            .O(N__22862),
            .I(N__22859));
    Odrv4 I__4552 (
            .O(N__22859),
            .I(\processor_zipi8.shift_rotate_result_7 ));
    InMux I__4551 (
            .O(N__22856),
            .I(N__22853));
    LocalMux I__4550 (
            .O(N__22853),
            .I(N__22850));
    Span4Mux_h I__4549 (
            .O(N__22850),
            .I(N__22847));
    Span4Mux_h I__4548 (
            .O(N__22847),
            .I(N__22844));
    Odrv4 I__4547 (
            .O(N__22844),
            .I(\processor_zipi8.spm_data_7 ));
    CascadeMux I__4546 (
            .O(N__22841),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269_cascade_ ));
    CascadeMux I__4545 (
            .O(N__22838),
            .I(N__22835));
    InMux I__4544 (
            .O(N__22835),
            .I(N__22829));
    InMux I__4543 (
            .O(N__22834),
            .I(N__22829));
    LocalMux I__4542 (
            .O(N__22829),
            .I(N__22826));
    Span4Mux_v I__4541 (
            .O(N__22826),
            .I(N__22823));
    Span4Mux_v I__4540 (
            .O(N__22823),
            .I(N__22820));
    Odrv4 I__4539 (
            .O(N__22820),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_7 ));
    InMux I__4538 (
            .O(N__22817),
            .I(N__22811));
    InMux I__4537 (
            .O(N__22816),
            .I(N__22811));
    LocalMux I__4536 (
            .O(N__22811),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_7 ));
    CascadeMux I__4535 (
            .O(N__22808),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_243_cascade_ ));
    InMux I__4534 (
            .O(N__22805),
            .I(N__22802));
    LocalMux I__4533 (
            .O(N__22802),
            .I(N__22799));
    Span4Mux_h I__4532 (
            .O(N__22799),
            .I(N__22796));
    Odrv4 I__4531 (
            .O(N__22796),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_299 ));
    CascadeMux I__4530 (
            .O(N__22793),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_5_cascade_ ));
    InMux I__4529 (
            .O(N__22790),
            .I(N__22787));
    LocalMux I__4528 (
            .O(N__22787),
            .I(N__22784));
    Span4Mux_s3_h I__4527 (
            .O(N__22784),
            .I(N__22781));
    Span4Mux_h I__4526 (
            .O(N__22781),
            .I(N__22778));
    Span4Mux_v I__4525 (
            .O(N__22778),
            .I(N__22775));
    Odrv4 I__4524 (
            .O(N__22775),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_315 ));
    InMux I__4523 (
            .O(N__22772),
            .I(N__22769));
    LocalMux I__4522 (
            .O(N__22769),
            .I(N__22765));
    InMux I__4521 (
            .O(N__22768),
            .I(N__22762));
    Span4Mux_v I__4520 (
            .O(N__22765),
            .I(N__22759));
    LocalMux I__4519 (
            .O(N__22762),
            .I(N__22756));
    Odrv4 I__4518 (
            .O(N__22759),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5 ));
    Odrv12 I__4517 (
            .O(N__22756),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5 ));
    CascadeMux I__4516 (
            .O(N__22751),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_5_cascade_ ));
    InMux I__4515 (
            .O(N__22748),
            .I(N__22744));
    InMux I__4514 (
            .O(N__22747),
            .I(N__22741));
    LocalMux I__4513 (
            .O(N__22744),
            .I(N__22736));
    LocalMux I__4512 (
            .O(N__22741),
            .I(N__22736));
    Span4Mux_v I__4511 (
            .O(N__22736),
            .I(N__22733));
    Odrv4 I__4510 (
            .O(N__22733),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_5 ));
    InMux I__4509 (
            .O(N__22730),
            .I(N__22727));
    LocalMux I__4508 (
            .O(N__22727),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_219 ));
    CascadeMux I__4507 (
            .O(N__22724),
            .I(N__22721));
    InMux I__4506 (
            .O(N__22721),
            .I(N__22718));
    LocalMux I__4505 (
            .O(N__22718),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_5 ));
    InMux I__4504 (
            .O(N__22715),
            .I(N__22712));
    LocalMux I__4503 (
            .O(N__22712),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_275 ));
    CascadeMux I__4502 (
            .O(N__22709),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_5_cascade_ ));
    InMux I__4501 (
            .O(N__22706),
            .I(N__22703));
    LocalMux I__4500 (
            .O(N__22703),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_5 ));
    CascadeMux I__4499 (
            .O(N__22700),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_5_cascade_ ));
    InMux I__4498 (
            .O(N__22697),
            .I(N__22694));
    LocalMux I__4497 (
            .O(N__22694),
            .I(N__22691));
    Span4Mux_v I__4496 (
            .O(N__22691),
            .I(N__22688));
    Span4Mux_h I__4495 (
            .O(N__22688),
            .I(N__22685));
    Odrv4 I__4494 (
            .O(N__22685),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_5 ));
    InMux I__4493 (
            .O(N__22682),
            .I(N__22679));
    LocalMux I__4492 (
            .O(N__22679),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_5 ));
    InMux I__4491 (
            .O(N__22676),
            .I(N__22673));
    LocalMux I__4490 (
            .O(N__22673),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_5 ));
    CascadeMux I__4489 (
            .O(N__22670),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_5_cascade_ ));
    InMux I__4488 (
            .O(N__22667),
            .I(N__22664));
    LocalMux I__4487 (
            .O(N__22664),
            .I(N__22660));
    InMux I__4486 (
            .O(N__22663),
            .I(N__22657));
    Odrv4 I__4485 (
            .O(N__22660),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5 ));
    LocalMux I__4484 (
            .O(N__22657),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5 ));
    InMux I__4483 (
            .O(N__22652),
            .I(N__22649));
    LocalMux I__4482 (
            .O(N__22649),
            .I(N__22645));
    InMux I__4481 (
            .O(N__22648),
            .I(N__22642));
    Span4Mux_h I__4480 (
            .O(N__22645),
            .I(N__22637));
    LocalMux I__4479 (
            .O(N__22642),
            .I(N__22637));
    Span4Mux_v I__4478 (
            .O(N__22637),
            .I(N__22634));
    Odrv4 I__4477 (
            .O(N__22634),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_5 ));
    CascadeMux I__4476 (
            .O(N__22631),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_5_cascade_ ));
    CascadeMux I__4475 (
            .O(N__22628),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_6_cascade_ ));
    InMux I__4474 (
            .O(N__22625),
            .I(N__22622));
    LocalMux I__4473 (
            .O(N__22622),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI0VUU1_6 ));
    CascadeMux I__4472 (
            .O(N__22619),
            .I(N__22616));
    InMux I__4471 (
            .O(N__22616),
            .I(N__22613));
    LocalMux I__4470 (
            .O(N__22613),
            .I(N__22610));
    Span4Mux_v I__4469 (
            .O(N__22610),
            .I(N__22606));
    InMux I__4468 (
            .O(N__22609),
            .I(N__22603));
    Odrv4 I__4467 (
            .O(N__22606),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6 ));
    LocalMux I__4466 (
            .O(N__22603),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6 ));
    InMux I__4465 (
            .O(N__22598),
            .I(N__22595));
    LocalMux I__4464 (
            .O(N__22595),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIQCIQ1_6 ));
    InMux I__4463 (
            .O(N__22592),
            .I(N__22588));
    InMux I__4462 (
            .O(N__22591),
            .I(N__22585));
    LocalMux I__4461 (
            .O(N__22588),
            .I(N__22582));
    LocalMux I__4460 (
            .O(N__22585),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6 ));
    Odrv4 I__4459 (
            .O(N__22582),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6 ));
    InMux I__4458 (
            .O(N__22577),
            .I(N__22571));
    InMux I__4457 (
            .O(N__22576),
            .I(N__22571));
    LocalMux I__4456 (
            .O(N__22571),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_7 ));
    SRMux I__4455 (
            .O(N__22568),
            .I(N__22564));
    SRMux I__4454 (
            .O(N__22567),
            .I(N__22557));
    LocalMux I__4453 (
            .O(N__22564),
            .I(N__22552));
    SRMux I__4452 (
            .O(N__22563),
            .I(N__22549));
    SRMux I__4451 (
            .O(N__22562),
            .I(N__22546));
    SRMux I__4450 (
            .O(N__22561),
            .I(N__22543));
    SRMux I__4449 (
            .O(N__22560),
            .I(N__22540));
    LocalMux I__4448 (
            .O(N__22557),
            .I(N__22537));
    SRMux I__4447 (
            .O(N__22556),
            .I(N__22534));
    SRMux I__4446 (
            .O(N__22555),
            .I(N__22531));
    Span4Mux_v I__4445 (
            .O(N__22552),
            .I(N__22524));
    LocalMux I__4444 (
            .O(N__22549),
            .I(N__22524));
    LocalMux I__4443 (
            .O(N__22546),
            .I(N__22521));
    LocalMux I__4442 (
            .O(N__22543),
            .I(N__22516));
    LocalMux I__4441 (
            .O(N__22540),
            .I(N__22516));
    Span4Mux_s2_v I__4440 (
            .O(N__22537),
            .I(N__22509));
    LocalMux I__4439 (
            .O(N__22534),
            .I(N__22509));
    LocalMux I__4438 (
            .O(N__22531),
            .I(N__22509));
    SRMux I__4437 (
            .O(N__22530),
            .I(N__22506));
    SRMux I__4436 (
            .O(N__22529),
            .I(N__22503));
    Span4Mux_v I__4435 (
            .O(N__22524),
            .I(N__22498));
    Span4Mux_v I__4434 (
            .O(N__22521),
            .I(N__22493));
    Span4Mux_v I__4433 (
            .O(N__22516),
            .I(N__22493));
    Span4Mux_v I__4432 (
            .O(N__22509),
            .I(N__22486));
    LocalMux I__4431 (
            .O(N__22506),
            .I(N__22486));
    LocalMux I__4430 (
            .O(N__22503),
            .I(N__22486));
    SRMux I__4429 (
            .O(N__22502),
            .I(N__22483));
    SRMux I__4428 (
            .O(N__22501),
            .I(N__22480));
    Span4Mux_v I__4427 (
            .O(N__22498),
            .I(N__22476));
    Span4Mux_v I__4426 (
            .O(N__22493),
            .I(N__22473));
    Span4Mux_v I__4425 (
            .O(N__22486),
            .I(N__22466));
    LocalMux I__4424 (
            .O(N__22483),
            .I(N__22466));
    LocalMux I__4423 (
            .O(N__22480),
            .I(N__22466));
    SRMux I__4422 (
            .O(N__22479),
            .I(N__22463));
    Sp12to4 I__4421 (
            .O(N__22476),
            .I(N__22460));
    Span4Mux_h I__4420 (
            .O(N__22473),
            .I(N__22457));
    Span4Mux_v I__4419 (
            .O(N__22466),
            .I(N__22454));
    LocalMux I__4418 (
            .O(N__22463),
            .I(N__22451));
    Odrv12 I__4417 (
            .O(N__22460),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4416 (
            .O(N__22457),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4415 (
            .O(N__22454),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4414 (
            .O(N__22451),
            .I(CONSTANT_ONE_NET));
    InMux I__4413 (
            .O(N__22442),
            .I(N__22439));
    LocalMux I__4412 (
            .O(N__22439),
            .I(N__22435));
    InMux I__4411 (
            .O(N__22438),
            .I(N__22432));
    Span4Mux_v I__4410 (
            .O(N__22435),
            .I(N__22429));
    LocalMux I__4409 (
            .O(N__22432),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6 ));
    Odrv4 I__4408 (
            .O(N__22429),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6 ));
    CascadeMux I__4407 (
            .O(N__22424),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_6_cascade_ ));
    CascadeMux I__4406 (
            .O(N__22421),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNICIK32_6_cascade_ ));
    CascadeMux I__4405 (
            .O(N__22418),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_6_cascade_ ));
    InMux I__4404 (
            .O(N__22415),
            .I(N__22412));
    LocalMux I__4403 (
            .O(N__22412),
            .I(N__22409));
    Span4Mux_h I__4402 (
            .O(N__22409),
            .I(N__22406));
    Odrv4 I__4401 (
            .O(N__22406),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFJCI8_6 ));
    InMux I__4400 (
            .O(N__22403),
            .I(N__22400));
    LocalMux I__4399 (
            .O(N__22400),
            .I(N__22396));
    InMux I__4398 (
            .O(N__22399),
            .I(N__22393));
    Odrv4 I__4397 (
            .O(N__22396),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2 ));
    LocalMux I__4396 (
            .O(N__22393),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2 ));
    InMux I__4395 (
            .O(N__22388),
            .I(N__22384));
    InMux I__4394 (
            .O(N__22387),
            .I(N__22381));
    LocalMux I__4393 (
            .O(N__22384),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3 ));
    LocalMux I__4392 (
            .O(N__22381),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3 ));
    InMux I__4391 (
            .O(N__22376),
            .I(N__22372));
    InMux I__4390 (
            .O(N__22375),
            .I(N__22369));
    LocalMux I__4389 (
            .O(N__22372),
            .I(N__22364));
    LocalMux I__4388 (
            .O(N__22369),
            .I(N__22364));
    Span4Mux_h I__4387 (
            .O(N__22364),
            .I(N__22361));
    Span4Mux_v I__4386 (
            .O(N__22361),
            .I(N__22358));
    Span4Mux_v I__4385 (
            .O(N__22358),
            .I(N__22355));
    Odrv4 I__4384 (
            .O(N__22355),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_6 ));
    CEMux I__4383 (
            .O(N__22352),
            .I(N__22349));
    LocalMux I__4382 (
            .O(N__22349),
            .I(N__22346));
    Span4Mux_s3_v I__4381 (
            .O(N__22346),
            .I(N__22343));
    Span4Mux_v I__4380 (
            .O(N__22343),
            .I(N__22340));
    Span4Mux_v I__4379 (
            .O(N__22340),
            .I(N__22336));
    CEMux I__4378 (
            .O(N__22339),
            .I(N__22333));
    Odrv4 I__4377 (
            .O(N__22336),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7 ));
    LocalMux I__4376 (
            .O(N__22333),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7 ));
    InMux I__4375 (
            .O(N__22328),
            .I(N__22325));
    LocalMux I__4374 (
            .O(N__22325),
            .I(N__22322));
    Span4Mux_h I__4373 (
            .O(N__22322),
            .I(N__22319));
    Span4Mux_v I__4372 (
            .O(N__22319),
            .I(N__22316));
    Odrv4 I__4371 (
            .O(N__22316),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI0ESR1_2 ));
    CascadeMux I__4370 (
            .O(N__22313),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_2_cascade_ ));
    InMux I__4369 (
            .O(N__22310),
            .I(N__22307));
    LocalMux I__4368 (
            .O(N__22307),
            .I(N__22304));
    Span4Mux_v I__4367 (
            .O(N__22304),
            .I(N__22301));
    Span4Mux_v I__4366 (
            .O(N__22301),
            .I(N__22298));
    Odrv4 I__4365 (
            .O(N__22298),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI2HMP1_2 ));
    CascadeMux I__4364 (
            .O(N__22295),
            .I(N__22280));
    CascadeMux I__4363 (
            .O(N__22294),
            .I(N__22276));
    CascadeMux I__4362 (
            .O(N__22293),
            .I(N__22273));
    CascadeMux I__4361 (
            .O(N__22292),
            .I(N__22269));
    CascadeMux I__4360 (
            .O(N__22291),
            .I(N__22263));
    CascadeMux I__4359 (
            .O(N__22290),
            .I(N__22259));
    CascadeMux I__4358 (
            .O(N__22289),
            .I(N__22256));
    CascadeMux I__4357 (
            .O(N__22288),
            .I(N__22252));
    CascadeMux I__4356 (
            .O(N__22287),
            .I(N__22248));
    CascadeMux I__4355 (
            .O(N__22286),
            .I(N__22242));
    CascadeMux I__4354 (
            .O(N__22285),
            .I(N__22238));
    CascadeMux I__4353 (
            .O(N__22284),
            .I(N__22235));
    CascadeMux I__4352 (
            .O(N__22283),
            .I(N__22227));
    InMux I__4351 (
            .O(N__22280),
            .I(N__22210));
    InMux I__4350 (
            .O(N__22279),
            .I(N__22210));
    InMux I__4349 (
            .O(N__22276),
            .I(N__22210));
    InMux I__4348 (
            .O(N__22273),
            .I(N__22210));
    InMux I__4347 (
            .O(N__22272),
            .I(N__22210));
    InMux I__4346 (
            .O(N__22269),
            .I(N__22210));
    InMux I__4345 (
            .O(N__22268),
            .I(N__22210));
    InMux I__4344 (
            .O(N__22267),
            .I(N__22210));
    InMux I__4343 (
            .O(N__22266),
            .I(N__22193));
    InMux I__4342 (
            .O(N__22263),
            .I(N__22193));
    InMux I__4341 (
            .O(N__22262),
            .I(N__22193));
    InMux I__4340 (
            .O(N__22259),
            .I(N__22193));
    InMux I__4339 (
            .O(N__22256),
            .I(N__22193));
    InMux I__4338 (
            .O(N__22255),
            .I(N__22193));
    InMux I__4337 (
            .O(N__22252),
            .I(N__22193));
    InMux I__4336 (
            .O(N__22251),
            .I(N__22193));
    InMux I__4335 (
            .O(N__22248),
            .I(N__22176));
    InMux I__4334 (
            .O(N__22247),
            .I(N__22176));
    InMux I__4333 (
            .O(N__22246),
            .I(N__22176));
    InMux I__4332 (
            .O(N__22245),
            .I(N__22176));
    InMux I__4331 (
            .O(N__22242),
            .I(N__22176));
    InMux I__4330 (
            .O(N__22241),
            .I(N__22176));
    InMux I__4329 (
            .O(N__22238),
            .I(N__22176));
    InMux I__4328 (
            .O(N__22235),
            .I(N__22176));
    InMux I__4327 (
            .O(N__22234),
            .I(N__22173));
    InMux I__4326 (
            .O(N__22233),
            .I(N__22170));
    InMux I__4325 (
            .O(N__22232),
            .I(N__22166));
    InMux I__4324 (
            .O(N__22231),
            .I(N__22163));
    InMux I__4323 (
            .O(N__22230),
            .I(N__22160));
    InMux I__4322 (
            .O(N__22227),
            .I(N__22156));
    LocalMux I__4321 (
            .O(N__22210),
            .I(N__22151));
    LocalMux I__4320 (
            .O(N__22193),
            .I(N__22151));
    LocalMux I__4319 (
            .O(N__22176),
            .I(N__22146));
    LocalMux I__4318 (
            .O(N__22173),
            .I(N__22146));
    LocalMux I__4317 (
            .O(N__22170),
            .I(N__22143));
    InMux I__4316 (
            .O(N__22169),
            .I(N__22140));
    LocalMux I__4315 (
            .O(N__22166),
            .I(N__22129));
    LocalMux I__4314 (
            .O(N__22163),
            .I(N__22124));
    LocalMux I__4313 (
            .O(N__22160),
            .I(N__22124));
    InMux I__4312 (
            .O(N__22159),
            .I(N__22121));
    LocalMux I__4311 (
            .O(N__22156),
            .I(N__22116));
    Sp12to4 I__4310 (
            .O(N__22151),
            .I(N__22116));
    Span4Mux_v I__4309 (
            .O(N__22146),
            .I(N__22113));
    Span4Mux_v I__4308 (
            .O(N__22143),
            .I(N__22110));
    LocalMux I__4307 (
            .O(N__22140),
            .I(N__22107));
    InMux I__4306 (
            .O(N__22139),
            .I(N__22092));
    InMux I__4305 (
            .O(N__22138),
            .I(N__22092));
    InMux I__4304 (
            .O(N__22137),
            .I(N__22092));
    InMux I__4303 (
            .O(N__22136),
            .I(N__22092));
    InMux I__4302 (
            .O(N__22135),
            .I(N__22092));
    InMux I__4301 (
            .O(N__22134),
            .I(N__22092));
    InMux I__4300 (
            .O(N__22133),
            .I(N__22092));
    InMux I__4299 (
            .O(N__22132),
            .I(N__22089));
    Span4Mux_s3_h I__4298 (
            .O(N__22129),
            .I(N__22082));
    Span4Mux_v I__4297 (
            .O(N__22124),
            .I(N__22082));
    LocalMux I__4296 (
            .O(N__22121),
            .I(N__22082));
    Span12Mux_v I__4295 (
            .O(N__22116),
            .I(N__22079));
    Span4Mux_v I__4294 (
            .O(N__22113),
            .I(N__22076));
    Span4Mux_v I__4293 (
            .O(N__22110),
            .I(N__22071));
    Span4Mux_s3_v I__4292 (
            .O(N__22107),
            .I(N__22071));
    LocalMux I__4291 (
            .O(N__22092),
            .I(N__22066));
    LocalMux I__4290 (
            .O(N__22089),
            .I(N__22066));
    Span4Mux_h I__4289 (
            .O(N__22082),
            .I(N__22063));
    Odrv12 I__4288 (
            .O(N__22079),
            .I(\processor_zipi8.sx_addr_4 ));
    Odrv4 I__4287 (
            .O(N__22076),
            .I(\processor_zipi8.sx_addr_4 ));
    Odrv4 I__4286 (
            .O(N__22071),
            .I(\processor_zipi8.sx_addr_4 ));
    Odrv12 I__4285 (
            .O(N__22066),
            .I(\processor_zipi8.sx_addr_4 ));
    Odrv4 I__4284 (
            .O(N__22063),
            .I(\processor_zipi8.sx_addr_4 ));
    CascadeMux I__4283 (
            .O(N__22052),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI792G8_2_cascade_ ));
    InMux I__4282 (
            .O(N__22049),
            .I(N__22046));
    LocalMux I__4281 (
            .O(N__22046),
            .I(N__22036));
    InMux I__4280 (
            .O(N__22045),
            .I(N__22031));
    InMux I__4279 (
            .O(N__22044),
            .I(N__22031));
    CascadeMux I__4278 (
            .O(N__22043),
            .I(N__22028));
    InMux I__4277 (
            .O(N__22042),
            .I(N__22019));
    InMux I__4276 (
            .O(N__22041),
            .I(N__22019));
    InMux I__4275 (
            .O(N__22040),
            .I(N__22019));
    InMux I__4274 (
            .O(N__22039),
            .I(N__22019));
    Span4Mux_s3_h I__4273 (
            .O(N__22036),
            .I(N__22014));
    LocalMux I__4272 (
            .O(N__22031),
            .I(N__22014));
    InMux I__4271 (
            .O(N__22028),
            .I(N__22010));
    LocalMux I__4270 (
            .O(N__22019),
            .I(N__22007));
    Span4Mux_v I__4269 (
            .O(N__22014),
            .I(N__22004));
    InMux I__4268 (
            .O(N__22013),
            .I(N__22001));
    LocalMux I__4267 (
            .O(N__22010),
            .I(N__21996));
    Span4Mux_h I__4266 (
            .O(N__22007),
            .I(N__21996));
    Span4Mux_h I__4265 (
            .O(N__22004),
            .I(N__21993));
    LocalMux I__4264 (
            .O(N__22001),
            .I(N__21990));
    Span4Mux_v I__4263 (
            .O(N__21996),
            .I(N__21987));
    Odrv4 I__4262 (
            .O(N__21993),
            .I(\processor_zipi8.sx_2 ));
    Odrv12 I__4261 (
            .O(N__21990),
            .I(\processor_zipi8.sx_2 ));
    Odrv4 I__4260 (
            .O(N__21987),
            .I(\processor_zipi8.sx_2 ));
    CascadeMux I__4259 (
            .O(N__21980),
            .I(N__21976));
    InMux I__4258 (
            .O(N__21979),
            .I(N__21973));
    InMux I__4257 (
            .O(N__21976),
            .I(N__21970));
    LocalMux I__4256 (
            .O(N__21973),
            .I(N__21965));
    LocalMux I__4255 (
            .O(N__21970),
            .I(N__21965));
    Odrv12 I__4254 (
            .O(N__21965),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_0 ));
    InMux I__4253 (
            .O(N__21962),
            .I(N__21959));
    LocalMux I__4252 (
            .O(N__21959),
            .I(N__21956));
    Span12Mux_s8_h I__4251 (
            .O(N__21956),
            .I(N__21953));
    Odrv12 I__4250 (
            .O(N__21953),
            .I(\processor_zipi8.shift_rotate_result_3 ));
    InMux I__4249 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__4248 (
            .O(N__21947),
            .I(N__21944));
    Span4Mux_h I__4247 (
            .O(N__21944),
            .I(N__21941));
    Span4Mux_v I__4246 (
            .O(N__21941),
            .I(N__21938));
    Odrv4 I__4245 (
            .O(N__21938),
            .I(\processor_zipi8.spm_data_3 ));
    CascadeMux I__4244 (
            .O(N__21935),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266_cascade_ ));
    InMux I__4243 (
            .O(N__21932),
            .I(N__21928));
    InMux I__4242 (
            .O(N__21931),
            .I(N__21925));
    LocalMux I__4241 (
            .O(N__21928),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3 ));
    LocalMux I__4240 (
            .O(N__21925),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3 ));
    CascadeMux I__4239 (
            .O(N__21920),
            .I(N__21917));
    InMux I__4238 (
            .O(N__21917),
            .I(N__21914));
    LocalMux I__4237 (
            .O(N__21914),
            .I(N__21910));
    InMux I__4236 (
            .O(N__21913),
            .I(N__21907));
    Span4Mux_v I__4235 (
            .O(N__21910),
            .I(N__21902));
    LocalMux I__4234 (
            .O(N__21907),
            .I(N__21902));
    Span4Mux_v I__4233 (
            .O(N__21902),
            .I(N__21899));
    Odrv4 I__4232 (
            .O(N__21899),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_0 ));
    InMux I__4231 (
            .O(N__21896),
            .I(N__21893));
    LocalMux I__4230 (
            .O(N__21893),
            .I(N__21890));
    Span4Mux_h I__4229 (
            .O(N__21890),
            .I(N__21887));
    Odrv4 I__4228 (
            .O(N__21887),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI8MSR1_4 ));
    CascadeMux I__4227 (
            .O(N__21884),
            .I(N__21881));
    InMux I__4226 (
            .O(N__21881),
            .I(N__21878));
    LocalMux I__4225 (
            .O(N__21878),
            .I(N__21875));
    Span4Mux_v I__4224 (
            .O(N__21875),
            .I(N__21872));
    Odrv4 I__4223 (
            .O(N__21872),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIAPMP1_4 ));
    InMux I__4222 (
            .O(N__21869),
            .I(N__21866));
    LocalMux I__4221 (
            .O(N__21866),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFIBI8_4 ));
    CascadeMux I__4220 (
            .O(N__21863),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7A3G8_4_cascade_ ));
    InMux I__4219 (
            .O(N__21860),
            .I(N__21857));
    LocalMux I__4218 (
            .O(N__21857),
            .I(N__21852));
    InMux I__4217 (
            .O(N__21856),
            .I(N__21847));
    InMux I__4216 (
            .O(N__21855),
            .I(N__21847));
    Span4Mux_v I__4215 (
            .O(N__21852),
            .I(N__21843));
    LocalMux I__4214 (
            .O(N__21847),
            .I(N__21840));
    InMux I__4213 (
            .O(N__21846),
            .I(N__21837));
    Span4Mux_s3_h I__4212 (
            .O(N__21843),
            .I(N__21828));
    Span4Mux_v I__4211 (
            .O(N__21840),
            .I(N__21828));
    LocalMux I__4210 (
            .O(N__21837),
            .I(N__21828));
    CascadeMux I__4209 (
            .O(N__21836),
            .I(N__21825));
    CascadeMux I__4208 (
            .O(N__21835),
            .I(N__21822));
    Span4Mux_h I__4207 (
            .O(N__21828),
            .I(N__21818));
    InMux I__4206 (
            .O(N__21825),
            .I(N__21811));
    InMux I__4205 (
            .O(N__21822),
            .I(N__21811));
    InMux I__4204 (
            .O(N__21821),
            .I(N__21811));
    Odrv4 I__4203 (
            .O(N__21818),
            .I(\processor_zipi8.sx_4 ));
    LocalMux I__4202 (
            .O(N__21811),
            .I(\processor_zipi8.sx_4 ));
    CascadeMux I__4201 (
            .O(N__21806),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNISRE42_4_cascade_ ));
    InMux I__4200 (
            .O(N__21803),
            .I(N__21800));
    LocalMux I__4199 (
            .O(N__21800),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_4 ));
    InMux I__4198 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__4197 (
            .O(N__21794),
            .I(N__21791));
    Span4Mux_v I__4196 (
            .O(N__21791),
            .I(N__21787));
    InMux I__4195 (
            .O(N__21790),
            .I(N__21784));
    Odrv4 I__4194 (
            .O(N__21787),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2 ));
    LocalMux I__4193 (
            .O(N__21784),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2 ));
    CascadeMux I__4192 (
            .O(N__21779),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_2_cascade_ ));
    CascadeMux I__4191 (
            .O(N__21776),
            .I(N__21773));
    InMux I__4190 (
            .O(N__21773),
            .I(N__21770));
    LocalMux I__4189 (
            .O(N__21770),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_2 ));
    InMux I__4188 (
            .O(N__21767),
            .I(N__21764));
    LocalMux I__4187 (
            .O(N__21764),
            .I(N__21761));
    Odrv4 I__4186 (
            .O(N__21761),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI4KGN1_2 ));
    CascadeMux I__4185 (
            .O(N__21758),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIKJE42_2_cascade_ ));
    CascadeMux I__4184 (
            .O(N__21755),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_1_cascade_ ));
    CascadeMux I__4183 (
            .O(N__21752),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_119_cascade_ ));
    CascadeMux I__4182 (
            .O(N__21749),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_1_cascade_ ));
    InMux I__4181 (
            .O(N__21746),
            .I(N__21743));
    LocalMux I__4180 (
            .O(N__21743),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_95 ));
    InMux I__4179 (
            .O(N__21740),
            .I(N__21737));
    LocalMux I__4178 (
            .O(N__21737),
            .I(N__21734));
    Odrv12 I__4177 (
            .O(N__21734),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_151 ));
    CascadeMux I__4176 (
            .O(N__21731),
            .I(N__21728));
    InMux I__4175 (
            .O(N__21728),
            .I(N__21725));
    LocalMux I__4174 (
            .O(N__21725),
            .I(N__21722));
    Span4Mux_h I__4173 (
            .O(N__21722),
            .I(N__21719));
    Odrv4 I__4172 (
            .O(N__21719),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_175 ));
    InMux I__4171 (
            .O(N__21716),
            .I(N__21713));
    LocalMux I__4170 (
            .O(N__21713),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_1 ));
    CascadeMux I__4169 (
            .O(N__21710),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_191_cascade_ ));
    InMux I__4168 (
            .O(N__21707),
            .I(N__21703));
    InMux I__4167 (
            .O(N__21706),
            .I(N__21698));
    LocalMux I__4166 (
            .O(N__21703),
            .I(N__21695));
    InMux I__4165 (
            .O(N__21702),
            .I(N__21690));
    InMux I__4164 (
            .O(N__21701),
            .I(N__21690));
    LocalMux I__4163 (
            .O(N__21698),
            .I(N__21687));
    Span4Mux_h I__4162 (
            .O(N__21695),
            .I(N__21677));
    LocalMux I__4161 (
            .O(N__21690),
            .I(N__21677));
    Span4Mux_v I__4160 (
            .O(N__21687),
            .I(N__21674));
    InMux I__4159 (
            .O(N__21686),
            .I(N__21669));
    InMux I__4158 (
            .O(N__21685),
            .I(N__21669));
    InMux I__4157 (
            .O(N__21684),
            .I(N__21662));
    InMux I__4156 (
            .O(N__21683),
            .I(N__21662));
    InMux I__4155 (
            .O(N__21682),
            .I(N__21662));
    Span4Mux_v I__4154 (
            .O(N__21677),
            .I(N__21655));
    Span4Mux_h I__4153 (
            .O(N__21674),
            .I(N__21655));
    LocalMux I__4152 (
            .O(N__21669),
            .I(N__21655));
    LocalMux I__4151 (
            .O(N__21662),
            .I(\processor_zipi8.sx_1 ));
    Odrv4 I__4150 (
            .O(N__21655),
            .I(\processor_zipi8.sx_1 ));
    CascadeMux I__4149 (
            .O(N__21650),
            .I(N__21647));
    InMux I__4148 (
            .O(N__21647),
            .I(N__21644));
    LocalMux I__4147 (
            .O(N__21644),
            .I(N__21641));
    Odrv12 I__4146 (
            .O(N__21641),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNII4IQ1_4 ));
    CascadeMux I__4145 (
            .O(N__21638),
            .I(N__21635));
    InMux I__4144 (
            .O(N__21635),
            .I(N__21632));
    LocalMux I__4143 (
            .O(N__21632),
            .I(N__21629));
    Span4Mux_h I__4142 (
            .O(N__21629),
            .I(N__21626));
    Odrv4 I__4141 (
            .O(N__21626),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_4 ));
    InMux I__4140 (
            .O(N__21623),
            .I(N__21620));
    LocalMux I__4139 (
            .O(N__21620),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI4AK32_4 ));
    CascadeMux I__4138 (
            .O(N__21617),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIOMUU1_4_cascade_ ));
    InMux I__4137 (
            .O(N__21614),
            .I(N__21611));
    LocalMux I__4136 (
            .O(N__21611),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_4 ));
    InMux I__4135 (
            .O(N__21608),
            .I(N__21604));
    InMux I__4134 (
            .O(N__21607),
            .I(N__21601));
    LocalMux I__4133 (
            .O(N__21604),
            .I(N__21598));
    LocalMux I__4132 (
            .O(N__21601),
            .I(N__21595));
    Span4Mux_v I__4131 (
            .O(N__21598),
            .I(N__21592));
    Odrv4 I__4130 (
            .O(N__21595),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7 ));
    Odrv4 I__4129 (
            .O(N__21592),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7 ));
    InMux I__4128 (
            .O(N__21587),
            .I(N__21584));
    LocalMux I__4127 (
            .O(N__21584),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_7 ));
    InMux I__4126 (
            .O(N__21581),
            .I(N__21575));
    InMux I__4125 (
            .O(N__21580),
            .I(N__21575));
    LocalMux I__4124 (
            .O(N__21575),
            .I(N__21572));
    Odrv12 I__4123 (
            .O(N__21572),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_7 ));
    CascadeMux I__4122 (
            .O(N__21569),
            .I(N__21566));
    InMux I__4121 (
            .O(N__21566),
            .I(N__21562));
    CascadeMux I__4120 (
            .O(N__21565),
            .I(N__21559));
    LocalMux I__4119 (
            .O(N__21562),
            .I(N__21556));
    InMux I__4118 (
            .O(N__21559),
            .I(N__21553));
    Span4Mux_v I__4117 (
            .O(N__21556),
            .I(N__21548));
    LocalMux I__4116 (
            .O(N__21553),
            .I(N__21548));
    Span4Mux_h I__4115 (
            .O(N__21548),
            .I(N__21543));
    InMux I__4114 (
            .O(N__21547),
            .I(N__21538));
    InMux I__4113 (
            .O(N__21546),
            .I(N__21538));
    Odrv4 I__4112 (
            .O(N__21543),
            .I(\processor_zipi8.port_id_1 ));
    LocalMux I__4111 (
            .O(N__21538),
            .I(\processor_zipi8.port_id_1 ));
    InMux I__4110 (
            .O(N__21533),
            .I(N__21530));
    LocalMux I__4109 (
            .O(N__21530),
            .I(N__21527));
    Span4Mux_h I__4108 (
            .O(N__21527),
            .I(N__21524));
    Span4Mux_h I__4107 (
            .O(N__21524),
            .I(N__21521));
    Odrv4 I__4106 (
            .O(N__21521),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_1 ));
    InMux I__4105 (
            .O(N__21518),
            .I(N__21509));
    InMux I__4104 (
            .O(N__21517),
            .I(N__21509));
    InMux I__4103 (
            .O(N__21516),
            .I(N__21509));
    LocalMux I__4102 (
            .O(N__21509),
            .I(N__21504));
    InMux I__4101 (
            .O(N__21508),
            .I(N__21499));
    InMux I__4100 (
            .O(N__21507),
            .I(N__21499));
    Span4Mux_h I__4099 (
            .O(N__21504),
            .I(N__21494));
    LocalMux I__4098 (
            .O(N__21499),
            .I(N__21494));
    Span4Mux_v I__4097 (
            .O(N__21494),
            .I(N__21491));
    Span4Mux_v I__4096 (
            .O(N__21491),
            .I(N__21488));
    Span4Mux_s1_v I__4095 (
            .O(N__21488),
            .I(N__21485));
    Odrv4 I__4094 (
            .O(N__21485),
            .I(instruction_1));
    InMux I__4093 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__4092 (
            .O(N__21479),
            .I(N__21476));
    Span4Mux_h I__4091 (
            .O(N__21476),
            .I(N__21473));
    Odrv4 I__4090 (
            .O(N__21473),
            .I(\processor_zipi8.pc_vector_1 ));
    InMux I__4089 (
            .O(N__21470),
            .I(N__21467));
    LocalMux I__4088 (
            .O(N__21467),
            .I(N__21464));
    Span4Mux_h I__4087 (
            .O(N__21464),
            .I(N__21461));
    Odrv4 I__4086 (
            .O(N__21461),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_4 ));
    CascadeMux I__4085 (
            .O(N__21458),
            .I(N__21449));
    CascadeMux I__4084 (
            .O(N__21457),
            .I(N__21433));
    InMux I__4083 (
            .O(N__21456),
            .I(N__21429));
    InMux I__4082 (
            .O(N__21455),
            .I(N__21424));
    InMux I__4081 (
            .O(N__21454),
            .I(N__21424));
    InMux I__4080 (
            .O(N__21453),
            .I(N__21421));
    InMux I__4079 (
            .O(N__21452),
            .I(N__21418));
    InMux I__4078 (
            .O(N__21449),
            .I(N__21411));
    InMux I__4077 (
            .O(N__21448),
            .I(N__21411));
    InMux I__4076 (
            .O(N__21447),
            .I(N__21406));
    InMux I__4075 (
            .O(N__21446),
            .I(N__21406));
    InMux I__4074 (
            .O(N__21445),
            .I(N__21403));
    InMux I__4073 (
            .O(N__21444),
            .I(N__21392));
    InMux I__4072 (
            .O(N__21443),
            .I(N__21392));
    InMux I__4071 (
            .O(N__21442),
            .I(N__21392));
    InMux I__4070 (
            .O(N__21441),
            .I(N__21383));
    InMux I__4069 (
            .O(N__21440),
            .I(N__21383));
    InMux I__4068 (
            .O(N__21439),
            .I(N__21380));
    InMux I__4067 (
            .O(N__21438),
            .I(N__21375));
    InMux I__4066 (
            .O(N__21437),
            .I(N__21375));
    InMux I__4065 (
            .O(N__21436),
            .I(N__21372));
    InMux I__4064 (
            .O(N__21433),
            .I(N__21369));
    InMux I__4063 (
            .O(N__21432),
            .I(N__21366));
    LocalMux I__4062 (
            .O(N__21429),
            .I(N__21357));
    LocalMux I__4061 (
            .O(N__21424),
            .I(N__21357));
    LocalMux I__4060 (
            .O(N__21421),
            .I(N__21357));
    LocalMux I__4059 (
            .O(N__21418),
            .I(N__21357));
    InMux I__4058 (
            .O(N__21417),
            .I(N__21350));
    InMux I__4057 (
            .O(N__21416),
            .I(N__21350));
    LocalMux I__4056 (
            .O(N__21411),
            .I(N__21345));
    LocalMux I__4055 (
            .O(N__21406),
            .I(N__21345));
    LocalMux I__4054 (
            .O(N__21403),
            .I(N__21342));
    InMux I__4053 (
            .O(N__21402),
            .I(N__21337));
    InMux I__4052 (
            .O(N__21401),
            .I(N__21337));
    InMux I__4051 (
            .O(N__21400),
            .I(N__21332));
    InMux I__4050 (
            .O(N__21399),
            .I(N__21332));
    LocalMux I__4049 (
            .O(N__21392),
            .I(N__21329));
    InMux I__4048 (
            .O(N__21391),
            .I(N__21326));
    InMux I__4047 (
            .O(N__21390),
            .I(N__21319));
    InMux I__4046 (
            .O(N__21389),
            .I(N__21319));
    InMux I__4045 (
            .O(N__21388),
            .I(N__21319));
    LocalMux I__4044 (
            .O(N__21383),
            .I(N__21316));
    LocalMux I__4043 (
            .O(N__21380),
            .I(N__21311));
    LocalMux I__4042 (
            .O(N__21375),
            .I(N__21311));
    LocalMux I__4041 (
            .O(N__21372),
            .I(N__21306));
    LocalMux I__4040 (
            .O(N__21369),
            .I(N__21306));
    LocalMux I__4039 (
            .O(N__21366),
            .I(N__21301));
    Span4Mux_v I__4038 (
            .O(N__21357),
            .I(N__21301));
    InMux I__4037 (
            .O(N__21356),
            .I(N__21296));
    InMux I__4036 (
            .O(N__21355),
            .I(N__21296));
    LocalMux I__4035 (
            .O(N__21350),
            .I(N__21293));
    Span4Mux_h I__4034 (
            .O(N__21345),
            .I(N__21284));
    Span4Mux_v I__4033 (
            .O(N__21342),
            .I(N__21284));
    LocalMux I__4032 (
            .O(N__21337),
            .I(N__21284));
    LocalMux I__4031 (
            .O(N__21332),
            .I(N__21284));
    Span4Mux_s3_v I__4030 (
            .O(N__21329),
            .I(N__21281));
    LocalMux I__4029 (
            .O(N__21326),
            .I(N__21274));
    LocalMux I__4028 (
            .O(N__21319),
            .I(N__21274));
    Span4Mux_h I__4027 (
            .O(N__21316),
            .I(N__21274));
    Span4Mux_s3_v I__4026 (
            .O(N__21311),
            .I(N__21271));
    Span4Mux_s3_v I__4025 (
            .O(N__21306),
            .I(N__21260));
    Span4Mux_h I__4024 (
            .O(N__21301),
            .I(N__21260));
    LocalMux I__4023 (
            .O(N__21296),
            .I(N__21260));
    Span4Mux_s3_v I__4022 (
            .O(N__21293),
            .I(N__21260));
    Span4Mux_v I__4021 (
            .O(N__21284),
            .I(N__21260));
    Span4Mux_h I__4020 (
            .O(N__21281),
            .I(N__21253));
    Span4Mux_v I__4019 (
            .O(N__21274),
            .I(N__21253));
    Span4Mux_h I__4018 (
            .O(N__21271),
            .I(N__21253));
    Span4Mux_h I__4017 (
            .O(N__21260),
            .I(N__21250));
    Odrv4 I__4016 (
            .O(N__21253),
            .I(instruction_12));
    Odrv4 I__4015 (
            .O(N__21250),
            .I(instruction_12));
    InMux I__4014 (
            .O(N__21245),
            .I(N__21239));
    InMux I__4013 (
            .O(N__21244),
            .I(N__21239));
    LocalMux I__4012 (
            .O(N__21239),
            .I(N__21236));
    Span4Mux_v I__4011 (
            .O(N__21236),
            .I(N__21233));
    Span4Mux_h I__4010 (
            .O(N__21233),
            .I(N__21230));
    Odrv4 I__4009 (
            .O(N__21230),
            .I(\processor_zipi8.pc_vector_4 ));
    InMux I__4008 (
            .O(N__21227),
            .I(N__21220));
    InMux I__4007 (
            .O(N__21226),
            .I(N__21217));
    InMux I__4006 (
            .O(N__21225),
            .I(N__21204));
    InMux I__4005 (
            .O(N__21224),
            .I(N__21204));
    InMux I__4004 (
            .O(N__21223),
            .I(N__21204));
    LocalMux I__4003 (
            .O(N__21220),
            .I(N__21201));
    LocalMux I__4002 (
            .O(N__21217),
            .I(N__21198));
    InMux I__4001 (
            .O(N__21216),
            .I(N__21193));
    InMux I__4000 (
            .O(N__21215),
            .I(N__21193));
    InMux I__3999 (
            .O(N__21214),
            .I(N__21190));
    CascadeMux I__3998 (
            .O(N__21213),
            .I(N__21186));
    CascadeMux I__3997 (
            .O(N__21212),
            .I(N__21183));
    InMux I__3996 (
            .O(N__21211),
            .I(N__21176));
    LocalMux I__3995 (
            .O(N__21204),
            .I(N__21171));
    Span4Mux_v I__3994 (
            .O(N__21201),
            .I(N__21171));
    Span4Mux_h I__3993 (
            .O(N__21198),
            .I(N__21164));
    LocalMux I__3992 (
            .O(N__21193),
            .I(N__21164));
    LocalMux I__3991 (
            .O(N__21190),
            .I(N__21164));
    InMux I__3990 (
            .O(N__21189),
            .I(N__21157));
    InMux I__3989 (
            .O(N__21186),
            .I(N__21157));
    InMux I__3988 (
            .O(N__21183),
            .I(N__21157));
    InMux I__3987 (
            .O(N__21182),
            .I(N__21152));
    InMux I__3986 (
            .O(N__21181),
            .I(N__21152));
    InMux I__3985 (
            .O(N__21180),
            .I(N__21147));
    InMux I__3984 (
            .O(N__21179),
            .I(N__21147));
    LocalMux I__3983 (
            .O(N__21176),
            .I(N__21144));
    Span4Mux_v I__3982 (
            .O(N__21171),
            .I(N__21135));
    Span4Mux_v I__3981 (
            .O(N__21164),
            .I(N__21135));
    LocalMux I__3980 (
            .O(N__21157),
            .I(N__21135));
    LocalMux I__3979 (
            .O(N__21152),
            .I(N__21135));
    LocalMux I__3978 (
            .O(N__21147),
            .I(N__21132));
    Span4Mux_s2_v I__3977 (
            .O(N__21144),
            .I(N__21129));
    Span4Mux_s2_v I__3976 (
            .O(N__21135),
            .I(N__21124));
    Span4Mux_h I__3975 (
            .O(N__21132),
            .I(N__21124));
    Span4Mux_h I__3974 (
            .O(N__21129),
            .I(N__21121));
    Span4Mux_h I__3973 (
            .O(N__21124),
            .I(N__21118));
    Odrv4 I__3972 (
            .O(N__21121),
            .I(instruction_13));
    Odrv4 I__3971 (
            .O(N__21118),
            .I(instruction_13));
    InMux I__3970 (
            .O(N__21113),
            .I(N__21107));
    InMux I__3969 (
            .O(N__21112),
            .I(N__21103));
    InMux I__3968 (
            .O(N__21111),
            .I(N__21100));
    InMux I__3967 (
            .O(N__21110),
            .I(N__21097));
    LocalMux I__3966 (
            .O(N__21107),
            .I(N__21094));
    InMux I__3965 (
            .O(N__21106),
            .I(N__21091));
    LocalMux I__3964 (
            .O(N__21103),
            .I(N__21087));
    LocalMux I__3963 (
            .O(N__21100),
            .I(N__21084));
    LocalMux I__3962 (
            .O(N__21097),
            .I(N__21075));
    Span4Mux_s3_h I__3961 (
            .O(N__21094),
            .I(N__21072));
    LocalMux I__3960 (
            .O(N__21091),
            .I(N__21069));
    InMux I__3959 (
            .O(N__21090),
            .I(N__21066));
    Span4Mux_v I__3958 (
            .O(N__21087),
            .I(N__21061));
    Span4Mux_s3_h I__3957 (
            .O(N__21084),
            .I(N__21061));
    InMux I__3956 (
            .O(N__21083),
            .I(N__21058));
    InMux I__3955 (
            .O(N__21082),
            .I(N__21047));
    InMux I__3954 (
            .O(N__21081),
            .I(N__21047));
    InMux I__3953 (
            .O(N__21080),
            .I(N__21047));
    InMux I__3952 (
            .O(N__21079),
            .I(N__21047));
    InMux I__3951 (
            .O(N__21078),
            .I(N__21047));
    Odrv12 I__3950 (
            .O(N__21075),
            .I(\processor_zipi8.sx_0 ));
    Odrv4 I__3949 (
            .O(N__21072),
            .I(\processor_zipi8.sx_0 ));
    Odrv4 I__3948 (
            .O(N__21069),
            .I(\processor_zipi8.sx_0 ));
    LocalMux I__3947 (
            .O(N__21066),
            .I(\processor_zipi8.sx_0 ));
    Odrv4 I__3946 (
            .O(N__21061),
            .I(\processor_zipi8.sx_0 ));
    LocalMux I__3945 (
            .O(N__21058),
            .I(\processor_zipi8.sx_0 ));
    LocalMux I__3944 (
            .O(N__21047),
            .I(\processor_zipi8.sx_0 ));
    IoInMux I__3943 (
            .O(N__21032),
            .I(N__21029));
    LocalMux I__3942 (
            .O(N__21029),
            .I(N__21026));
    IoSpan4Mux I__3941 (
            .O(N__21026),
            .I(N__21023));
    Span4Mux_s3_h I__3940 (
            .O(N__21023),
            .I(N__21020));
    Odrv4 I__3939 (
            .O(N__21020),
            .I(LED1_c));
    InMux I__3938 (
            .O(N__21017),
            .I(N__21011));
    InMux I__3937 (
            .O(N__21016),
            .I(N__21011));
    LocalMux I__3936 (
            .O(N__21011),
            .I(N__21008));
    Span12Mux_s10_h I__3935 (
            .O(N__21008),
            .I(N__21005));
    Odrv12 I__3934 (
            .O(N__21005),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_1 ));
    CascadeMux I__3933 (
            .O(N__21002),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_1_cascade_ ));
    InMux I__3932 (
            .O(N__20999),
            .I(N__20993));
    InMux I__3931 (
            .O(N__20998),
            .I(N__20993));
    LocalMux I__3930 (
            .O(N__20993),
            .I(N__20990));
    Odrv12 I__3929 (
            .O(N__20990),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_1 ));
    InMux I__3928 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__3927 (
            .O(N__20984),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1 ));
    InMux I__3926 (
            .O(N__20981),
            .I(N__20975));
    InMux I__3925 (
            .O(N__20980),
            .I(N__20975));
    LocalMux I__3924 (
            .O(N__20975),
            .I(N__20972));
    Odrv4 I__3923 (
            .O(N__20972),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_1 ));
    CascadeMux I__3922 (
            .O(N__20969),
            .I(N__20966));
    InMux I__3921 (
            .O(N__20966),
            .I(N__20960));
    InMux I__3920 (
            .O(N__20965),
            .I(N__20960));
    LocalMux I__3919 (
            .O(N__20960),
            .I(N__20957));
    Span4Mux_v I__3918 (
            .O(N__20957),
            .I(N__20954));
    Odrv4 I__3917 (
            .O(N__20954),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_1 ));
    CascadeMux I__3916 (
            .O(N__20951),
            .I(N__20948));
    InMux I__3915 (
            .O(N__20948),
            .I(N__20945));
    LocalMux I__3914 (
            .O(N__20945),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_1 ));
    InMux I__3913 (
            .O(N__20942),
            .I(N__20939));
    LocalMux I__3912 (
            .O(N__20939),
            .I(N__20936));
    Odrv12 I__3911 (
            .O(N__20936),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_7 ));
    InMux I__3910 (
            .O(N__20933),
            .I(N__20930));
    LocalMux I__3909 (
            .O(N__20930),
            .I(N__20927));
    Span4Mux_s3_h I__3908 (
            .O(N__20927),
            .I(N__20924));
    Span4Mux_h I__3907 (
            .O(N__20924),
            .I(N__20921));
    Odrv4 I__3906 (
            .O(N__20921),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_7 ));
    CascadeMux I__3905 (
            .O(N__20918),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_0_cascade_ ));
    CascadeMux I__3904 (
            .O(N__20915),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_0_cascade_ ));
    CascadeMux I__3903 (
            .O(N__20912),
            .I(N__20909));
    InMux I__3902 (
            .O(N__20909),
            .I(N__20906));
    LocalMux I__3901 (
            .O(N__20906),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_7 ));
    CascadeMux I__3900 (
            .O(N__20903),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_0_cascade_ ));
    InMux I__3899 (
            .O(N__20900),
            .I(N__20897));
    LocalMux I__3898 (
            .O(N__20897),
            .I(N__20893));
    InMux I__3897 (
            .O(N__20896),
            .I(N__20890));
    Span4Mux_v I__3896 (
            .O(N__20893),
            .I(N__20885));
    LocalMux I__3895 (
            .O(N__20890),
            .I(N__20885));
    Span4Mux_v I__3894 (
            .O(N__20885),
            .I(N__20882));
    Odrv4 I__3893 (
            .O(N__20882),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_0 ));
    InMux I__3892 (
            .O(N__20879),
            .I(N__20876));
    LocalMux I__3891 (
            .O(N__20876),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_0 ));
    InMux I__3890 (
            .O(N__20873),
            .I(N__20867));
    InMux I__3889 (
            .O(N__20872),
            .I(N__20867));
    LocalMux I__3888 (
            .O(N__20867),
            .I(N__20864));
    Span4Mux_h I__3887 (
            .O(N__20864),
            .I(N__20861));
    Odrv4 I__3886 (
            .O(N__20861),
            .I(\processor_zipi8.register_enable ));
    CascadeMux I__3885 (
            .O(N__20858),
            .I(N__20843));
    InMux I__3884 (
            .O(N__20857),
            .I(N__20832));
    InMux I__3883 (
            .O(N__20856),
            .I(N__20832));
    InMux I__3882 (
            .O(N__20855),
            .I(N__20832));
    InMux I__3881 (
            .O(N__20854),
            .I(N__20832));
    InMux I__3880 (
            .O(N__20853),
            .I(N__20828));
    InMux I__3879 (
            .O(N__20852),
            .I(N__20813));
    InMux I__3878 (
            .O(N__20851),
            .I(N__20813));
    InMux I__3877 (
            .O(N__20850),
            .I(N__20813));
    InMux I__3876 (
            .O(N__20849),
            .I(N__20813));
    InMux I__3875 (
            .O(N__20848),
            .I(N__20813));
    InMux I__3874 (
            .O(N__20847),
            .I(N__20813));
    InMux I__3873 (
            .O(N__20846),
            .I(N__20813));
    InMux I__3872 (
            .O(N__20843),
            .I(N__20808));
    InMux I__3871 (
            .O(N__20842),
            .I(N__20808));
    InMux I__3870 (
            .O(N__20841),
            .I(N__20805));
    LocalMux I__3869 (
            .O(N__20832),
            .I(N__20802));
    InMux I__3868 (
            .O(N__20831),
            .I(N__20799));
    LocalMux I__3867 (
            .O(N__20828),
            .I(N__20794));
    LocalMux I__3866 (
            .O(N__20813),
            .I(N__20794));
    LocalMux I__3865 (
            .O(N__20808),
            .I(N__20787));
    LocalMux I__3864 (
            .O(N__20805),
            .I(N__20787));
    Span4Mux_v I__3863 (
            .O(N__20802),
            .I(N__20787));
    LocalMux I__3862 (
            .O(N__20799),
            .I(N__20782));
    Sp12to4 I__3861 (
            .O(N__20794),
            .I(N__20782));
    Odrv4 I__3860 (
            .O(N__20787),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205 ));
    Odrv12 I__3859 (
            .O(N__20782),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205 ));
    InMux I__3858 (
            .O(N__20777),
            .I(N__20774));
    LocalMux I__3857 (
            .O(N__20774),
            .I(N__20771));
    Odrv4 I__3856 (
            .O(N__20771),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_0 ));
    InMux I__3855 (
            .O(N__20768),
            .I(N__20765));
    LocalMux I__3854 (
            .O(N__20765),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNISBGN1_0 ));
    CascadeMux I__3853 (
            .O(N__20762),
            .I(N__20759));
    InMux I__3852 (
            .O(N__20759),
            .I(N__20756));
    LocalMux I__3851 (
            .O(N__20756),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_1 ));
    InMux I__3850 (
            .O(N__20753),
            .I(N__20749));
    InMux I__3849 (
            .O(N__20752),
            .I(N__20746));
    LocalMux I__3848 (
            .O(N__20749),
            .I(N__20743));
    LocalMux I__3847 (
            .O(N__20746),
            .I(N__20740));
    Span4Mux_v I__3846 (
            .O(N__20743),
            .I(N__20735));
    Span4Mux_h I__3845 (
            .O(N__20740),
            .I(N__20735));
    Odrv4 I__3844 (
            .O(N__20735),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_1 ));
    InMux I__3843 (
            .O(N__20732),
            .I(N__20728));
    InMux I__3842 (
            .O(N__20731),
            .I(N__20725));
    LocalMux I__3841 (
            .O(N__20728),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1 ));
    LocalMux I__3840 (
            .O(N__20725),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1 ));
    CascadeMux I__3839 (
            .O(N__20720),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_1_cascade_ ));
    CascadeMux I__3838 (
            .O(N__20717),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_cascade_ ));
    InMux I__3837 (
            .O(N__20714),
            .I(N__20708));
    InMux I__3836 (
            .O(N__20713),
            .I(N__20708));
    LocalMux I__3835 (
            .O(N__20708),
            .I(N__20705));
    Span4Mux_v I__3834 (
            .O(N__20705),
            .I(N__20702));
    Span4Mux_h I__3833 (
            .O(N__20702),
            .I(N__20699));
    Odrv4 I__3832 (
            .O(N__20699),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_1 ));
    CascadeMux I__3831 (
            .O(N__20696),
            .I(N__20692));
    CascadeMux I__3830 (
            .O(N__20695),
            .I(N__20689));
    InMux I__3829 (
            .O(N__20692),
            .I(N__20684));
    InMux I__3828 (
            .O(N__20689),
            .I(N__20684));
    LocalMux I__3827 (
            .O(N__20684),
            .I(N__20681));
    Span4Mux_h I__3826 (
            .O(N__20681),
            .I(N__20678));
    Odrv4 I__3825 (
            .O(N__20678),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_1 ));
    InMux I__3824 (
            .O(N__20675),
            .I(N__20672));
    LocalMux I__3823 (
            .O(N__20672),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_5 ));
    CascadeMux I__3822 (
            .O(N__20669),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_5_cascade_ ));
    InMux I__3821 (
            .O(N__20666),
            .I(N__20663));
    LocalMux I__3820 (
            .O(N__20663),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_5 ));
    InMux I__3819 (
            .O(N__20660),
            .I(N__20648));
    InMux I__3818 (
            .O(N__20659),
            .I(N__20648));
    InMux I__3817 (
            .O(N__20658),
            .I(N__20648));
    InMux I__3816 (
            .O(N__20657),
            .I(N__20648));
    LocalMux I__3815 (
            .O(N__20648),
            .I(N__20635));
    CascadeMux I__3814 (
            .O(N__20647),
            .I(N__20632));
    CascadeMux I__3813 (
            .O(N__20646),
            .I(N__20629));
    InMux I__3812 (
            .O(N__20645),
            .I(N__20624));
    InMux I__3811 (
            .O(N__20644),
            .I(N__20609));
    InMux I__3810 (
            .O(N__20643),
            .I(N__20609));
    InMux I__3809 (
            .O(N__20642),
            .I(N__20609));
    InMux I__3808 (
            .O(N__20641),
            .I(N__20609));
    InMux I__3807 (
            .O(N__20640),
            .I(N__20609));
    InMux I__3806 (
            .O(N__20639),
            .I(N__20609));
    InMux I__3805 (
            .O(N__20638),
            .I(N__20609));
    Span4Mux_v I__3804 (
            .O(N__20635),
            .I(N__20606));
    InMux I__3803 (
            .O(N__20632),
            .I(N__20597));
    InMux I__3802 (
            .O(N__20629),
            .I(N__20597));
    InMux I__3801 (
            .O(N__20628),
            .I(N__20597));
    InMux I__3800 (
            .O(N__20627),
            .I(N__20597));
    LocalMux I__3799 (
            .O(N__20624),
            .I(N__20592));
    LocalMux I__3798 (
            .O(N__20609),
            .I(N__20592));
    Sp12to4 I__3797 (
            .O(N__20606),
            .I(N__20587));
    LocalMux I__3796 (
            .O(N__20597),
            .I(N__20587));
    Odrv4 I__3795 (
            .O(N__20592),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206 ));
    Odrv12 I__3794 (
            .O(N__20587),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206 ));
    CascadeMux I__3793 (
            .O(N__20582),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_0_cascade_ ));
    CascadeMux I__3792 (
            .O(N__20579),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNICBE42_0_cascade_ ));
    InMux I__3791 (
            .O(N__20576),
            .I(N__20573));
    LocalMux I__3790 (
            .O(N__20573),
            .I(N__20570));
    Span4Mux_v I__3789 (
            .O(N__20570),
            .I(N__20567));
    Odrv4 I__3788 (
            .O(N__20567),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIQ8MP1_0 ));
    CascadeMux I__3787 (
            .O(N__20564),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_0_cascade_ ));
    InMux I__3786 (
            .O(N__20561),
            .I(N__20558));
    LocalMux I__3785 (
            .O(N__20558),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIO5SR1_0 ));
    InMux I__3784 (
            .O(N__20555),
            .I(N__20552));
    LocalMux I__3783 (
            .O(N__20552),
            .I(N__20549));
    Span4Mux_h I__3782 (
            .O(N__20549),
            .I(N__20546));
    Odrv4 I__3781 (
            .O(N__20546),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI781G8_0 ));
    CascadeMux I__3780 (
            .O(N__20543),
            .I(N__20536));
    CascadeMux I__3779 (
            .O(N__20542),
            .I(N__20531));
    CascadeMux I__3778 (
            .O(N__20541),
            .I(N__20528));
    InMux I__3777 (
            .O(N__20540),
            .I(N__20524));
    InMux I__3776 (
            .O(N__20539),
            .I(N__20519));
    InMux I__3775 (
            .O(N__20536),
            .I(N__20519));
    InMux I__3774 (
            .O(N__20535),
            .I(N__20514));
    InMux I__3773 (
            .O(N__20534),
            .I(N__20514));
    InMux I__3772 (
            .O(N__20531),
            .I(N__20507));
    InMux I__3771 (
            .O(N__20528),
            .I(N__20507));
    InMux I__3770 (
            .O(N__20527),
            .I(N__20507));
    LocalMux I__3769 (
            .O(N__20524),
            .I(N__20502));
    LocalMux I__3768 (
            .O(N__20519),
            .I(N__20502));
    LocalMux I__3767 (
            .O(N__20514),
            .I(N__20497));
    LocalMux I__3766 (
            .O(N__20507),
            .I(N__20497));
    Span4Mux_v I__3765 (
            .O(N__20502),
            .I(N__20494));
    Odrv4 I__3764 (
            .O(N__20497),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209 ));
    Odrv4 I__3763 (
            .O(N__20494),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209 ));
    InMux I__3762 (
            .O(N__20489),
            .I(N__20486));
    LocalMux I__3761 (
            .O(N__20486),
            .I(N__20482));
    InMux I__3760 (
            .O(N__20485),
            .I(N__20479));
    Span4Mux_h I__3759 (
            .O(N__20482),
            .I(N__20474));
    LocalMux I__3758 (
            .O(N__20479),
            .I(N__20474));
    Span4Mux_v I__3757 (
            .O(N__20474),
            .I(N__20471));
    Odrv4 I__3756 (
            .O(N__20471),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_7 ));
    InMux I__3755 (
            .O(N__20468),
            .I(N__20462));
    InMux I__3754 (
            .O(N__20467),
            .I(N__20462));
    LocalMux I__3753 (
            .O(N__20462),
            .I(N__20459));
    Span4Mux_v I__3752 (
            .O(N__20459),
            .I(N__20456));
    Odrv4 I__3751 (
            .O(N__20456),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_7 ));
    InMux I__3750 (
            .O(N__20453),
            .I(N__20450));
    LocalMux I__3749 (
            .O(N__20450),
            .I(N__20447));
    Span4Mux_s3_h I__3748 (
            .O(N__20447),
            .I(N__20444));
    Odrv4 I__3747 (
            .O(N__20444),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_7 ));
    CascadeMux I__3746 (
            .O(N__20441),
            .I(N__20437));
    InMux I__3745 (
            .O(N__20440),
            .I(N__20432));
    InMux I__3744 (
            .O(N__20437),
            .I(N__20432));
    LocalMux I__3743 (
            .O(N__20432),
            .I(N__20429));
    Odrv4 I__3742 (
            .O(N__20429),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_7 ));
    InMux I__3741 (
            .O(N__20426),
            .I(N__20420));
    InMux I__3740 (
            .O(N__20425),
            .I(N__20420));
    LocalMux I__3739 (
            .O(N__20420),
            .I(N__20417));
    Span4Mux_v I__3738 (
            .O(N__20417),
            .I(N__20414));
    Odrv4 I__3737 (
            .O(N__20414),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_7 ));
    InMux I__3736 (
            .O(N__20411),
            .I(N__20408));
    LocalMux I__3735 (
            .O(N__20408),
            .I(N__20405));
    Odrv12 I__3734 (
            .O(N__20405),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_7 ));
    CascadeMux I__3733 (
            .O(N__20402),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_5_cascade_ ));
    InMux I__3732 (
            .O(N__20399),
            .I(N__20396));
    LocalMux I__3731 (
            .O(N__20396),
            .I(N__20393));
    Span12Mux_s6_h I__3730 (
            .O(N__20393),
            .I(N__20390));
    Odrv12 I__3729 (
            .O(N__20390),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_5 ));
    InMux I__3728 (
            .O(N__20387),
            .I(N__20383));
    InMux I__3727 (
            .O(N__20386),
            .I(N__20380));
    LocalMux I__3726 (
            .O(N__20383),
            .I(N__20377));
    LocalMux I__3725 (
            .O(N__20380),
            .I(N__20372));
    Span4Mux_v I__3724 (
            .O(N__20377),
            .I(N__20372));
    Odrv4 I__3723 (
            .O(N__20372),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_0 ));
    InMux I__3722 (
            .O(N__20369),
            .I(N__20365));
    InMux I__3721 (
            .O(N__20368),
            .I(N__20362));
    LocalMux I__3720 (
            .O(N__20365),
            .I(N__20359));
    LocalMux I__3719 (
            .O(N__20362),
            .I(N__20356));
    Span4Mux_h I__3718 (
            .O(N__20359),
            .I(N__20351));
    Span4Mux_v I__3717 (
            .O(N__20356),
            .I(N__20351));
    Odrv4 I__3716 (
            .O(N__20351),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_0 ));
    CascadeMux I__3715 (
            .O(N__20348),
            .I(N__20345));
    InMux I__3714 (
            .O(N__20345),
            .I(N__20342));
    LocalMux I__3713 (
            .O(N__20342),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_0 ));
    InMux I__3712 (
            .O(N__20339),
            .I(N__20336));
    LocalMux I__3711 (
            .O(N__20336),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_5 ));
    InMux I__3710 (
            .O(N__20333),
            .I(N__20327));
    InMux I__3709 (
            .O(N__20332),
            .I(N__20327));
    LocalMux I__3708 (
            .O(N__20327),
            .I(N__20321));
    CascadeMux I__3707 (
            .O(N__20326),
            .I(N__20318));
    CascadeMux I__3706 (
            .O(N__20325),
            .I(N__20313));
    CascadeMux I__3705 (
            .O(N__20324),
            .I(N__20310));
    Span4Mux_h I__3704 (
            .O(N__20321),
            .I(N__20307));
    InMux I__3703 (
            .O(N__20318),
            .I(N__20304));
    InMux I__3702 (
            .O(N__20317),
            .I(N__20295));
    InMux I__3701 (
            .O(N__20316),
            .I(N__20295));
    InMux I__3700 (
            .O(N__20313),
            .I(N__20295));
    InMux I__3699 (
            .O(N__20310),
            .I(N__20295));
    Odrv4 I__3698 (
            .O(N__20307),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212 ));
    LocalMux I__3697 (
            .O(N__20304),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212 ));
    LocalMux I__3696 (
            .O(N__20295),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212 ));
    CEMux I__3695 (
            .O(N__20288),
            .I(N__20284));
    CEMux I__3694 (
            .O(N__20287),
            .I(N__20281));
    LocalMux I__3693 (
            .O(N__20284),
            .I(N__20278));
    LocalMux I__3692 (
            .O(N__20281),
            .I(N__20275));
    Span4Mux_v I__3691 (
            .O(N__20278),
            .I(N__20272));
    Span4Mux_v I__3690 (
            .O(N__20275),
            .I(N__20269));
    Span4Mux_h I__3689 (
            .O(N__20272),
            .I(N__20266));
    Span4Mux_h I__3688 (
            .O(N__20269),
            .I(N__20263));
    Odrv4 I__3687 (
            .O(N__20266),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14 ));
    Odrv4 I__3686 (
            .O(N__20263),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14 ));
    CascadeMux I__3685 (
            .O(N__20258),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_4_cascade_ ));
    CascadeMux I__3684 (
            .O(N__20255),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_7_cascade_ ));
    CascadeMux I__3683 (
            .O(N__20252),
            .I(N__20249));
    InMux I__3682 (
            .O(N__20249),
            .I(N__20246));
    LocalMux I__3681 (
            .O(N__20246),
            .I(N__20243));
    Span12Mux_s6_h I__3680 (
            .O(N__20243),
            .I(N__20240));
    Odrv12 I__3679 (
            .O(N__20240),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIO8HN1_7 ));
    CascadeMux I__3678 (
            .O(N__20237),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_7_cascade_ ));
    CascadeMux I__3677 (
            .O(N__20234),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_7_cascade_ ));
    InMux I__3676 (
            .O(N__20231),
            .I(N__20228));
    LocalMux I__3675 (
            .O(N__20228),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI43VU1_7 ));
    CascadeMux I__3674 (
            .O(N__20225),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIGMK32_7_cascade_ ));
    InMux I__3673 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__3672 (
            .O(N__20219),
            .I(N__20216));
    Span4Mux_v I__3671 (
            .O(N__20216),
            .I(N__20213));
    Span4Mux_h I__3670 (
            .O(N__20213),
            .I(N__20210));
    Span4Mux_v I__3669 (
            .O(N__20210),
            .I(N__20207));
    Odrv4 I__3668 (
            .O(N__20207),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_7 ));
    InMux I__3667 (
            .O(N__20204),
            .I(N__20200));
    InMux I__3666 (
            .O(N__20203),
            .I(N__20197));
    LocalMux I__3665 (
            .O(N__20200),
            .I(N__20194));
    LocalMux I__3664 (
            .O(N__20197),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7 ));
    Odrv4 I__3663 (
            .O(N__20194),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7 ));
    CascadeMux I__3662 (
            .O(N__20189),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_7_cascade_ ));
    InMux I__3661 (
            .O(N__20186),
            .I(N__20180));
    InMux I__3660 (
            .O(N__20185),
            .I(N__20180));
    LocalMux I__3659 (
            .O(N__20180),
            .I(N__20177));
    Span4Mux_h I__3658 (
            .O(N__20177),
            .I(N__20174));
    Odrv4 I__3657 (
            .O(N__20174),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_7 ));
    InMux I__3656 (
            .O(N__20171),
            .I(N__20168));
    LocalMux I__3655 (
            .O(N__20168),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_7 ));
    InMux I__3654 (
            .O(N__20165),
            .I(N__20161));
    InMux I__3653 (
            .O(N__20164),
            .I(N__20158));
    LocalMux I__3652 (
            .O(N__20161),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3 ));
    LocalMux I__3651 (
            .O(N__20158),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3 ));
    CascadeMux I__3650 (
            .O(N__20153),
            .I(N__20150));
    InMux I__3649 (
            .O(N__20150),
            .I(N__20147));
    LocalMux I__3648 (
            .O(N__20147),
            .I(N__20144));
    Odrv4 I__3647 (
            .O(N__20144),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_3 ));
    CEMux I__3646 (
            .O(N__20141),
            .I(N__20137));
    CEMux I__3645 (
            .O(N__20140),
            .I(N__20134));
    LocalMux I__3644 (
            .O(N__20137),
            .I(N__20131));
    LocalMux I__3643 (
            .O(N__20134),
            .I(N__20128));
    Span4Mux_h I__3642 (
            .O(N__20131),
            .I(N__20125));
    Span4Mux_v I__3641 (
            .O(N__20128),
            .I(N__20122));
    Span4Mux_s1_v I__3640 (
            .O(N__20125),
            .I(N__20119));
    Span4Mux_v I__3639 (
            .O(N__20122),
            .I(N__20116));
    Odrv4 I__3638 (
            .O(N__20119),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6 ));
    Odrv4 I__3637 (
            .O(N__20116),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6 ));
    InMux I__3636 (
            .O(N__20111),
            .I(N__20108));
    LocalMux I__3635 (
            .O(N__20108),
            .I(\processor_zipi8.alu_result_4 ));
    CascadeMux I__3634 (
            .O(N__20105),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI8OGN1_3_cascade_ ));
    CascadeMux I__3633 (
            .O(N__20102),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_am_1_3_cascade_ ));
    InMux I__3632 (
            .O(N__20099),
            .I(N__20096));
    LocalMux I__3631 (
            .O(N__20096),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIONE42_3 ));
    InMux I__3630 (
            .O(N__20093),
            .I(N__20090));
    LocalMux I__3629 (
            .O(N__20090),
            .I(N__20087));
    Span12Mux_s3_v I__3628 (
            .O(N__20087),
            .I(N__20084));
    Odrv12 I__3627 (
            .O(N__20084),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI6LMP1_3 ));
    CascadeMux I__3626 (
            .O(N__20081),
            .I(N__20078));
    InMux I__3625 (
            .O(N__20078),
            .I(N__20075));
    LocalMux I__3624 (
            .O(N__20075),
            .I(N__20072));
    Span12Mux_s5_v I__3623 (
            .O(N__20072),
            .I(N__20069));
    Odrv12 I__3622 (
            .O(N__20069),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI4ISR1_3 ));
    InMux I__3621 (
            .O(N__20066),
            .I(N__20063));
    LocalMux I__3620 (
            .O(N__20063),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_3 ));
    CascadeMux I__3619 (
            .O(N__20060),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINP2G8_3_cascade_ ));
    CascadeMux I__3618 (
            .O(N__20057),
            .I(N__20053));
    InMux I__3617 (
            .O(N__20056),
            .I(N__20047));
    InMux I__3616 (
            .O(N__20053),
            .I(N__20040));
    InMux I__3615 (
            .O(N__20052),
            .I(N__20040));
    InMux I__3614 (
            .O(N__20051),
            .I(N__20037));
    InMux I__3613 (
            .O(N__20050),
            .I(N__20034));
    LocalMux I__3612 (
            .O(N__20047),
            .I(N__20031));
    CascadeMux I__3611 (
            .O(N__20046),
            .I(N__20028));
    CascadeMux I__3610 (
            .O(N__20045),
            .I(N__20025));
    LocalMux I__3609 (
            .O(N__20040),
            .I(N__20021));
    LocalMux I__3608 (
            .O(N__20037),
            .I(N__20018));
    LocalMux I__3607 (
            .O(N__20034),
            .I(N__20015));
    Span4Mux_h I__3606 (
            .O(N__20031),
            .I(N__20011));
    InMux I__3605 (
            .O(N__20028),
            .I(N__20004));
    InMux I__3604 (
            .O(N__20025),
            .I(N__20004));
    InMux I__3603 (
            .O(N__20024),
            .I(N__20004));
    Span12Mux_s5_h I__3602 (
            .O(N__20021),
            .I(N__20001));
    Span4Mux_h I__3601 (
            .O(N__20018),
            .I(N__19996));
    Span4Mux_v I__3600 (
            .O(N__20015),
            .I(N__19996));
    InMux I__3599 (
            .O(N__20014),
            .I(N__19993));
    Span4Mux_v I__3598 (
            .O(N__20011),
            .I(N__19988));
    LocalMux I__3597 (
            .O(N__20004),
            .I(N__19988));
    Odrv12 I__3596 (
            .O(N__20001),
            .I(\processor_zipi8.sx_3 ));
    Odrv4 I__3595 (
            .O(N__19996),
            .I(\processor_zipi8.sx_3 ));
    LocalMux I__3594 (
            .O(N__19993),
            .I(\processor_zipi8.sx_3 ));
    Odrv4 I__3593 (
            .O(N__19988),
            .I(\processor_zipi8.sx_3 ));
    InMux I__3592 (
            .O(N__19979),
            .I(N__19976));
    LocalMux I__3591 (
            .O(N__19976),
            .I(N__19973));
    Odrv12 I__3590 (
            .O(N__19973),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_4 ));
    InMux I__3589 (
            .O(N__19970),
            .I(N__19967));
    LocalMux I__3588 (
            .O(N__19967),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_4 ));
    CascadeMux I__3587 (
            .O(N__19964),
            .I(N__19960));
    InMux I__3586 (
            .O(N__19963),
            .I(N__19955));
    InMux I__3585 (
            .O(N__19960),
            .I(N__19952));
    CascadeMux I__3584 (
            .O(N__19959),
            .I(N__19940));
    CascadeMux I__3583 (
            .O(N__19958),
            .I(N__19933));
    LocalMux I__3582 (
            .O(N__19955),
            .I(N__19926));
    LocalMux I__3581 (
            .O(N__19952),
            .I(N__19926));
    InMux I__3580 (
            .O(N__19951),
            .I(N__19919));
    InMux I__3579 (
            .O(N__19950),
            .I(N__19919));
    InMux I__3578 (
            .O(N__19949),
            .I(N__19919));
    InMux I__3577 (
            .O(N__19948),
            .I(N__19914));
    InMux I__3576 (
            .O(N__19947),
            .I(N__19909));
    InMux I__3575 (
            .O(N__19946),
            .I(N__19909));
    InMux I__3574 (
            .O(N__19945),
            .I(N__19904));
    InMux I__3573 (
            .O(N__19944),
            .I(N__19904));
    InMux I__3572 (
            .O(N__19943),
            .I(N__19898));
    InMux I__3571 (
            .O(N__19940),
            .I(N__19887));
    InMux I__3570 (
            .O(N__19939),
            .I(N__19887));
    InMux I__3569 (
            .O(N__19938),
            .I(N__19887));
    InMux I__3568 (
            .O(N__19937),
            .I(N__19887));
    InMux I__3567 (
            .O(N__19936),
            .I(N__19887));
    InMux I__3566 (
            .O(N__19933),
            .I(N__19880));
    InMux I__3565 (
            .O(N__19932),
            .I(N__19880));
    InMux I__3564 (
            .O(N__19931),
            .I(N__19880));
    Span4Mux_v I__3563 (
            .O(N__19926),
            .I(N__19875));
    LocalMux I__3562 (
            .O(N__19919),
            .I(N__19875));
    InMux I__3561 (
            .O(N__19918),
            .I(N__19872));
    CascadeMux I__3560 (
            .O(N__19917),
            .I(N__19866));
    LocalMux I__3559 (
            .O(N__19914),
            .I(N__19859));
    LocalMux I__3558 (
            .O(N__19909),
            .I(N__19859));
    LocalMux I__3557 (
            .O(N__19904),
            .I(N__19859));
    InMux I__3556 (
            .O(N__19903),
            .I(N__19852));
    InMux I__3555 (
            .O(N__19902),
            .I(N__19852));
    InMux I__3554 (
            .O(N__19901),
            .I(N__19852));
    LocalMux I__3553 (
            .O(N__19898),
            .I(N__19845));
    LocalMux I__3552 (
            .O(N__19887),
            .I(N__19845));
    LocalMux I__3551 (
            .O(N__19880),
            .I(N__19845));
    Span4Mux_h I__3550 (
            .O(N__19875),
            .I(N__19842));
    LocalMux I__3549 (
            .O(N__19872),
            .I(N__19839));
    InMux I__3548 (
            .O(N__19871),
            .I(N__19830));
    InMux I__3547 (
            .O(N__19870),
            .I(N__19830));
    InMux I__3546 (
            .O(N__19869),
            .I(N__19830));
    InMux I__3545 (
            .O(N__19866),
            .I(N__19830));
    Span4Mux_v I__3544 (
            .O(N__19859),
            .I(N__19827));
    LocalMux I__3543 (
            .O(N__19852),
            .I(N__19824));
    Span4Mux_h I__3542 (
            .O(N__19845),
            .I(N__19819));
    Span4Mux_v I__3541 (
            .O(N__19842),
            .I(N__19819));
    Span4Mux_v I__3540 (
            .O(N__19839),
            .I(N__19816));
    LocalMux I__3539 (
            .O(N__19830),
            .I(N__19809));
    Sp12to4 I__3538 (
            .O(N__19827),
            .I(N__19809));
    Span12Mux_s2_h I__3537 (
            .O(N__19824),
            .I(N__19809));
    Span4Mux_h I__3536 (
            .O(N__19819),
            .I(N__19806));
    Odrv4 I__3535 (
            .O(N__19816),
            .I(instruction_14));
    Odrv12 I__3534 (
            .O(N__19809),
            .I(instruction_14));
    Odrv4 I__3533 (
            .O(N__19806),
            .I(instruction_14));
    InMux I__3532 (
            .O(N__19799),
            .I(N__19791));
    InMux I__3531 (
            .O(N__19798),
            .I(N__19788));
    InMux I__3530 (
            .O(N__19797),
            .I(N__19785));
    InMux I__3529 (
            .O(N__19796),
            .I(N__19771));
    InMux I__3528 (
            .O(N__19795),
            .I(N__19771));
    InMux I__3527 (
            .O(N__19794),
            .I(N__19768));
    LocalMux I__3526 (
            .O(N__19791),
            .I(N__19761));
    LocalMux I__3525 (
            .O(N__19788),
            .I(N__19761));
    LocalMux I__3524 (
            .O(N__19785),
            .I(N__19761));
    InMux I__3523 (
            .O(N__19784),
            .I(N__19758));
    InMux I__3522 (
            .O(N__19783),
            .I(N__19755));
    CascadeMux I__3521 (
            .O(N__19782),
            .I(N__19752));
    InMux I__3520 (
            .O(N__19781),
            .I(N__19744));
    InMux I__3519 (
            .O(N__19780),
            .I(N__19744));
    InMux I__3518 (
            .O(N__19779),
            .I(N__19744));
    CascadeMux I__3517 (
            .O(N__19778),
            .I(N__19740));
    InMux I__3516 (
            .O(N__19777),
            .I(N__19734));
    InMux I__3515 (
            .O(N__19776),
            .I(N__19734));
    LocalMux I__3514 (
            .O(N__19771),
            .I(N__19729));
    LocalMux I__3513 (
            .O(N__19768),
            .I(N__19729));
    Span4Mux_v I__3512 (
            .O(N__19761),
            .I(N__19722));
    LocalMux I__3511 (
            .O(N__19758),
            .I(N__19722));
    LocalMux I__3510 (
            .O(N__19755),
            .I(N__19722));
    InMux I__3509 (
            .O(N__19752),
            .I(N__19717));
    InMux I__3508 (
            .O(N__19751),
            .I(N__19717));
    LocalMux I__3507 (
            .O(N__19744),
            .I(N__19714));
    InMux I__3506 (
            .O(N__19743),
            .I(N__19709));
    InMux I__3505 (
            .O(N__19740),
            .I(N__19709));
    InMux I__3504 (
            .O(N__19739),
            .I(N__19706));
    LocalMux I__3503 (
            .O(N__19734),
            .I(N__19701));
    Span4Mux_h I__3502 (
            .O(N__19729),
            .I(N__19701));
    Span4Mux_h I__3501 (
            .O(N__19722),
            .I(N__19698));
    LocalMux I__3500 (
            .O(N__19717),
            .I(N__19691));
    Span4Mux_h I__3499 (
            .O(N__19714),
            .I(N__19691));
    LocalMux I__3498 (
            .O(N__19709),
            .I(N__19691));
    LocalMux I__3497 (
            .O(N__19706),
            .I(\processor_zipi8.arith_logical_sel_1_0_2 ));
    Odrv4 I__3496 (
            .O(N__19701),
            .I(\processor_zipi8.arith_logical_sel_1_0_2 ));
    Odrv4 I__3495 (
            .O(N__19698),
            .I(\processor_zipi8.arith_logical_sel_1_0_2 ));
    Odrv4 I__3494 (
            .O(N__19691),
            .I(\processor_zipi8.arith_logical_sel_1_0_2 ));
    InMux I__3493 (
            .O(N__19682),
            .I(N__19679));
    LocalMux I__3492 (
            .O(N__19679),
            .I(N__19676));
    Span12Mux_s6_v I__3491 (
            .O(N__19676),
            .I(N__19673));
    Odrv12 I__3490 (
            .O(N__19673),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_3 ));
    CascadeMux I__3489 (
            .O(N__19670),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_3_cascade_ ));
    CascadeMux I__3488 (
            .O(N__19667),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_3_cascade_ ));
    InMux I__3487 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__3486 (
            .O(N__19661),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_3 ));
    InMux I__3485 (
            .O(N__19658),
            .I(N__19655));
    LocalMux I__3484 (
            .O(N__19655),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_3 ));
    InMux I__3483 (
            .O(N__19652),
            .I(N__19646));
    InMux I__3482 (
            .O(N__19651),
            .I(N__19646));
    LocalMux I__3481 (
            .O(N__19646),
            .I(\processor_zipi8.sy_3 ));
    CascadeMux I__3480 (
            .O(N__19643),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_bm_1_3_cascade_ ));
    InMux I__3479 (
            .O(N__19640),
            .I(N__19636));
    InMux I__3478 (
            .O(N__19639),
            .I(N__19633));
    LocalMux I__3477 (
            .O(N__19636),
            .I(N__19628));
    LocalMux I__3476 (
            .O(N__19633),
            .I(N__19625));
    InMux I__3475 (
            .O(N__19632),
            .I(N__19622));
    InMux I__3474 (
            .O(N__19631),
            .I(N__19619));
    Span4Mux_v I__3473 (
            .O(N__19628),
            .I(N__19614));
    Span12Mux_s9_v I__3472 (
            .O(N__19625),
            .I(N__19609));
    LocalMux I__3471 (
            .O(N__19622),
            .I(N__19609));
    LocalMux I__3470 (
            .O(N__19619),
            .I(N__19606));
    InMux I__3469 (
            .O(N__19618),
            .I(N__19603));
    InMux I__3468 (
            .O(N__19617),
            .I(N__19600));
    Odrv4 I__3467 (
            .O(N__19614),
            .I(\processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical ));
    Odrv12 I__3466 (
            .O(N__19609),
            .I(\processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical ));
    Odrv12 I__3465 (
            .O(N__19606),
            .I(\processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical ));
    LocalMux I__3464 (
            .O(N__19603),
            .I(\processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical ));
    LocalMux I__3463 (
            .O(N__19600),
            .I(\processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical ));
    InMux I__3462 (
            .O(N__19589),
            .I(N__19581));
    InMux I__3461 (
            .O(N__19588),
            .I(N__19581));
    InMux I__3460 (
            .O(N__19587),
            .I(N__19572));
    InMux I__3459 (
            .O(N__19586),
            .I(N__19572));
    LocalMux I__3458 (
            .O(N__19581),
            .I(N__19569));
    InMux I__3457 (
            .O(N__19580),
            .I(N__19564));
    InMux I__3456 (
            .O(N__19579),
            .I(N__19564));
    InMux I__3455 (
            .O(N__19578),
            .I(N__19558));
    InMux I__3454 (
            .O(N__19577),
            .I(N__19558));
    LocalMux I__3453 (
            .O(N__19572),
            .I(N__19552));
    Span4Mux_v I__3452 (
            .O(N__19569),
            .I(N__19546));
    LocalMux I__3451 (
            .O(N__19564),
            .I(N__19546));
    InMux I__3450 (
            .O(N__19563),
            .I(N__19543));
    LocalMux I__3449 (
            .O(N__19558),
            .I(N__19540));
    InMux I__3448 (
            .O(N__19557),
            .I(N__19537));
    CascadeMux I__3447 (
            .O(N__19556),
            .I(N__19533));
    CascadeMux I__3446 (
            .O(N__19555),
            .I(N__19530));
    Span4Mux_v I__3445 (
            .O(N__19552),
            .I(N__19527));
    InMux I__3444 (
            .O(N__19551),
            .I(N__19524));
    Span4Mux_h I__3443 (
            .O(N__19546),
            .I(N__19515));
    LocalMux I__3442 (
            .O(N__19543),
            .I(N__19515));
    Span4Mux_v I__3441 (
            .O(N__19540),
            .I(N__19515));
    LocalMux I__3440 (
            .O(N__19537),
            .I(N__19515));
    InMux I__3439 (
            .O(N__19536),
            .I(N__19508));
    InMux I__3438 (
            .O(N__19533),
            .I(N__19508));
    InMux I__3437 (
            .O(N__19530),
            .I(N__19508));
    Odrv4 I__3436 (
            .O(N__19527),
            .I(\processor_zipi8.un4_arith_logical_sel ));
    LocalMux I__3435 (
            .O(N__19524),
            .I(\processor_zipi8.un4_arith_logical_sel ));
    Odrv4 I__3434 (
            .O(N__19515),
            .I(\processor_zipi8.un4_arith_logical_sel ));
    LocalMux I__3433 (
            .O(N__19508),
            .I(\processor_zipi8.un4_arith_logical_sel ));
    InMux I__3432 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__3431 (
            .O(N__19496),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1Z0Z_1 ));
    InMux I__3430 (
            .O(N__19493),
            .I(N__19490));
    LocalMux I__3429 (
            .O(N__19490),
            .I(\processor_zipi8.arith_and_logic_operations_i.N_773_tz ));
    CascadeMux I__3428 (
            .O(N__19487),
            .I(N__19483));
    InMux I__3427 (
            .O(N__19486),
            .I(N__19479));
    InMux I__3426 (
            .O(N__19483),
            .I(N__19475));
    CascadeMux I__3425 (
            .O(N__19482),
            .I(N__19468));
    LocalMux I__3424 (
            .O(N__19479),
            .I(N__19464));
    InMux I__3423 (
            .O(N__19478),
            .I(N__19461));
    LocalMux I__3422 (
            .O(N__19475),
            .I(N__19458));
    InMux I__3421 (
            .O(N__19474),
            .I(N__19454));
    InMux I__3420 (
            .O(N__19473),
            .I(N__19451));
    InMux I__3419 (
            .O(N__19472),
            .I(N__19444));
    InMux I__3418 (
            .O(N__19471),
            .I(N__19444));
    InMux I__3417 (
            .O(N__19468),
            .I(N__19444));
    InMux I__3416 (
            .O(N__19467),
            .I(N__19441));
    Span4Mux_v I__3415 (
            .O(N__19464),
            .I(N__19434));
    LocalMux I__3414 (
            .O(N__19461),
            .I(N__19434));
    Span4Mux_v I__3413 (
            .O(N__19458),
            .I(N__19434));
    InMux I__3412 (
            .O(N__19457),
            .I(N__19431));
    LocalMux I__3411 (
            .O(N__19454),
            .I(N__19428));
    LocalMux I__3410 (
            .O(N__19451),
            .I(N__19425));
    LocalMux I__3409 (
            .O(N__19444),
            .I(N__19420));
    LocalMux I__3408 (
            .O(N__19441),
            .I(N__19420));
    Span4Mux_h I__3407 (
            .O(N__19434),
            .I(N__19415));
    LocalMux I__3406 (
            .O(N__19431),
            .I(N__19415));
    Span12Mux_v I__3405 (
            .O(N__19428),
            .I(N__19412));
    Span4Mux_v I__3404 (
            .O(N__19425),
            .I(N__19407));
    Span4Mux_v I__3403 (
            .O(N__19420),
            .I(N__19407));
    Span4Mux_v I__3402 (
            .O(N__19415),
            .I(N__19404));
    Odrv12 I__3401 (
            .O(N__19412),
            .I(\processor_zipi8.arith_logical_sel_1_0_0 ));
    Odrv4 I__3400 (
            .O(N__19407),
            .I(\processor_zipi8.arith_logical_sel_1_0_0 ));
    Odrv4 I__3399 (
            .O(N__19404),
            .I(\processor_zipi8.arith_logical_sel_1_0_0 ));
    InMux I__3398 (
            .O(N__19397),
            .I(N__19394));
    LocalMux I__3397 (
            .O(N__19394),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_1 ));
    CascadeMux I__3396 (
            .O(N__19391),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_4_cascade_ ));
    InMux I__3395 (
            .O(N__19388),
            .I(N__19385));
    LocalMux I__3394 (
            .O(N__19385),
            .I(N__19382));
    Odrv4 I__3393 (
            .O(N__19382),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_4 ));
    CascadeMux I__3392 (
            .O(N__19379),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_4_cascade_ ));
    InMux I__3391 (
            .O(N__19376),
            .I(N__19370));
    InMux I__3390 (
            .O(N__19375),
            .I(N__19370));
    LocalMux I__3389 (
            .O(N__19370),
            .I(N__19367));
    Span4Mux_v I__3388 (
            .O(N__19367),
            .I(N__19364));
    Span4Mux_v I__3387 (
            .O(N__19364),
            .I(N__19361));
    Odrv4 I__3386 (
            .O(N__19361),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_4 ));
    InMux I__3385 (
            .O(N__19358),
            .I(N__19355));
    LocalMux I__3384 (
            .O(N__19355),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_4 ));
    InMux I__3383 (
            .O(N__19352),
            .I(N__19349));
    LocalMux I__3382 (
            .O(N__19349),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_4 ));
    CascadeMux I__3381 (
            .O(N__19346),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_4_cascade_ ));
    InMux I__3380 (
            .O(N__19343),
            .I(N__19340));
    LocalMux I__3379 (
            .O(N__19340),
            .I(N__19337));
    Odrv4 I__3378 (
            .O(N__19337),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_4 ));
    CascadeMux I__3377 (
            .O(N__19334),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4_cascade_ ));
    InMux I__3376 (
            .O(N__19331),
            .I(N__19325));
    InMux I__3375 (
            .O(N__19330),
            .I(N__19325));
    LocalMux I__3374 (
            .O(N__19325),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_34_5 ));
    InMux I__3373 (
            .O(N__19322),
            .I(N__19316));
    InMux I__3372 (
            .O(N__19321),
            .I(N__19316));
    LocalMux I__3371 (
            .O(N__19316),
            .I(N__19313));
    Odrv12 I__3370 (
            .O(N__19313),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_5 ));
    InMux I__3369 (
            .O(N__19310),
            .I(N__19307));
    LocalMux I__3368 (
            .O(N__19307),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4 ));
    InMux I__3367 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__3366 (
            .O(N__19301),
            .I(\processor_zipi8.flags_i.parity_5 ));
    CascadeMux I__3365 (
            .O(N__19298),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_1_cascade_ ));
    InMux I__3364 (
            .O(N__19295),
            .I(N__19291));
    InMux I__3363 (
            .O(N__19294),
            .I(N__19288));
    LocalMux I__3362 (
            .O(N__19291),
            .I(\processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1 ));
    LocalMux I__3361 (
            .O(N__19288),
            .I(\processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1 ));
    InMux I__3360 (
            .O(N__19283),
            .I(N__19280));
    LocalMux I__3359 (
            .O(N__19280),
            .I(N__19276));
    InMux I__3358 (
            .O(N__19279),
            .I(N__19273));
    Odrv12 I__3357 (
            .O(N__19276),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1 ));
    LocalMux I__3356 (
            .O(N__19273),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1 ));
    InMux I__3355 (
            .O(N__19268),
            .I(N__19265));
    LocalMux I__3354 (
            .O(N__19265),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tzZ0Z_4 ));
    CascadeMux I__3353 (
            .O(N__19262),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_4_cascade_ ));
    CascadeMux I__3352 (
            .O(N__19259),
            .I(N__19255));
    InMux I__3351 (
            .O(N__19258),
            .I(N__19250));
    InMux I__3350 (
            .O(N__19255),
            .I(N__19250));
    LocalMux I__3349 (
            .O(N__19250),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_4 ));
    CascadeMux I__3348 (
            .O(N__19247),
            .I(N__19243));
    CascadeMux I__3347 (
            .O(N__19246),
            .I(N__19240));
    InMux I__3346 (
            .O(N__19243),
            .I(N__19237));
    InMux I__3345 (
            .O(N__19240),
            .I(N__19231));
    LocalMux I__3344 (
            .O(N__19237),
            .I(N__19228));
    InMux I__3343 (
            .O(N__19236),
            .I(N__19221));
    InMux I__3342 (
            .O(N__19235),
            .I(N__19221));
    InMux I__3341 (
            .O(N__19234),
            .I(N__19221));
    LocalMux I__3340 (
            .O(N__19231),
            .I(N__19218));
    Span4Mux_h I__3339 (
            .O(N__19228),
            .I(N__19213));
    LocalMux I__3338 (
            .O(N__19221),
            .I(N__19213));
    Odrv4 I__3337 (
            .O(N__19218),
            .I(\processor_zipi8.port_id_4 ));
    Odrv4 I__3336 (
            .O(N__19213),
            .I(\processor_zipi8.port_id_4 ));
    InMux I__3335 (
            .O(N__19208),
            .I(N__19195));
    InMux I__3334 (
            .O(N__19207),
            .I(N__19195));
    InMux I__3333 (
            .O(N__19206),
            .I(N__19190));
    InMux I__3332 (
            .O(N__19205),
            .I(N__19190));
    InMux I__3331 (
            .O(N__19204),
            .I(N__19181));
    InMux I__3330 (
            .O(N__19203),
            .I(N__19181));
    CascadeMux I__3329 (
            .O(N__19202),
            .I(N__19177));
    InMux I__3328 (
            .O(N__19201),
            .I(N__19172));
    InMux I__3327 (
            .O(N__19200),
            .I(N__19172));
    LocalMux I__3326 (
            .O(N__19195),
            .I(N__19167));
    LocalMux I__3325 (
            .O(N__19190),
            .I(N__19167));
    InMux I__3324 (
            .O(N__19189),
            .I(N__19160));
    InMux I__3323 (
            .O(N__19188),
            .I(N__19160));
    InMux I__3322 (
            .O(N__19187),
            .I(N__19160));
    InMux I__3321 (
            .O(N__19186),
            .I(N__19157));
    LocalMux I__3320 (
            .O(N__19181),
            .I(N__19154));
    InMux I__3319 (
            .O(N__19180),
            .I(N__19147));
    InMux I__3318 (
            .O(N__19177),
            .I(N__19147));
    LocalMux I__3317 (
            .O(N__19172),
            .I(N__19144));
    Span4Mux_h I__3316 (
            .O(N__19167),
            .I(N__19137));
    LocalMux I__3315 (
            .O(N__19160),
            .I(N__19137));
    LocalMux I__3314 (
            .O(N__19157),
            .I(N__19137));
    Span4Mux_v I__3313 (
            .O(N__19154),
            .I(N__19134));
    InMux I__3312 (
            .O(N__19153),
            .I(N__19129));
    InMux I__3311 (
            .O(N__19152),
            .I(N__19129));
    LocalMux I__3310 (
            .O(N__19147),
            .I(N__19126));
    Span4Mux_v I__3309 (
            .O(N__19144),
            .I(N__19121));
    Span4Mux_v I__3308 (
            .O(N__19137),
            .I(N__19121));
    Odrv4 I__3307 (
            .O(N__19134),
            .I(\processor_zipi8.arith_logical_sel_1 ));
    LocalMux I__3306 (
            .O(N__19129),
            .I(\processor_zipi8.arith_logical_sel_1 ));
    Odrv12 I__3305 (
            .O(N__19126),
            .I(\processor_zipi8.arith_logical_sel_1 ));
    Odrv4 I__3304 (
            .O(N__19121),
            .I(\processor_zipi8.arith_logical_sel_1 ));
    InMux I__3303 (
            .O(N__19112),
            .I(N__19109));
    LocalMux I__3302 (
            .O(N__19109),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_4 ));
    CascadeMux I__3301 (
            .O(N__19106),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198_cascade_ ));
    InMux I__3300 (
            .O(N__19103),
            .I(N__19099));
    InMux I__3299 (
            .O(N__19102),
            .I(N__19096));
    LocalMux I__3298 (
            .O(N__19099),
            .I(N__19093));
    LocalMux I__3297 (
            .O(N__19096),
            .I(N__19090));
    Odrv4 I__3296 (
            .O(N__19093),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3 ));
    Odrv4 I__3295 (
            .O(N__19090),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3 ));
    InMux I__3294 (
            .O(N__19085),
            .I(N__19082));
    LocalMux I__3293 (
            .O(N__19082),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2 ));
    CascadeMux I__3292 (
            .O(N__19079),
            .I(N__19076));
    InMux I__3291 (
            .O(N__19076),
            .I(N__19073));
    LocalMux I__3290 (
            .O(N__19073),
            .I(\processor_zipi8.decode4_strobes_enables_i.un8_register_enable_type ));
    CEMux I__3289 (
            .O(N__19070),
            .I(N__19062));
    CascadeMux I__3288 (
            .O(N__19069),
            .I(N__19053));
    InMux I__3287 (
            .O(N__19068),
            .I(N__19046));
    InMux I__3286 (
            .O(N__19067),
            .I(N__19046));
    InMux I__3285 (
            .O(N__19066),
            .I(N__19046));
    InMux I__3284 (
            .O(N__19065),
            .I(N__19043));
    LocalMux I__3283 (
            .O(N__19062),
            .I(N__19038));
    InMux I__3282 (
            .O(N__19061),
            .I(N__19035));
    InMux I__3281 (
            .O(N__19060),
            .I(N__19032));
    CascadeMux I__3280 (
            .O(N__19059),
            .I(N__19028));
    InMux I__3279 (
            .O(N__19058),
            .I(N__19025));
    InMux I__3278 (
            .O(N__19057),
            .I(N__19018));
    InMux I__3277 (
            .O(N__19056),
            .I(N__19018));
    InMux I__3276 (
            .O(N__19053),
            .I(N__19018));
    LocalMux I__3275 (
            .O(N__19046),
            .I(N__19013));
    LocalMux I__3274 (
            .O(N__19043),
            .I(N__19013));
    InMux I__3273 (
            .O(N__19042),
            .I(N__19010));
    CascadeMux I__3272 (
            .O(N__19041),
            .I(N__19006));
    Span4Mux_v I__3271 (
            .O(N__19038),
            .I(N__19002));
    LocalMux I__3270 (
            .O(N__19035),
            .I(N__18995));
    LocalMux I__3269 (
            .O(N__19032),
            .I(N__18995));
    InMux I__3268 (
            .O(N__19031),
            .I(N__18992));
    InMux I__3267 (
            .O(N__19028),
            .I(N__18989));
    LocalMux I__3266 (
            .O(N__19025),
            .I(N__18980));
    LocalMux I__3265 (
            .O(N__19018),
            .I(N__18980));
    Span4Mux_h I__3264 (
            .O(N__19013),
            .I(N__18980));
    LocalMux I__3263 (
            .O(N__19010),
            .I(N__18980));
    InMux I__3262 (
            .O(N__19009),
            .I(N__18977));
    InMux I__3261 (
            .O(N__19006),
            .I(N__18972));
    InMux I__3260 (
            .O(N__19005),
            .I(N__18972));
    Span4Mux_s2_h I__3259 (
            .O(N__19002),
            .I(N__18969));
    InMux I__3258 (
            .O(N__19001),
            .I(N__18964));
    InMux I__3257 (
            .O(N__19000),
            .I(N__18964));
    Span4Mux_v I__3256 (
            .O(N__18995),
            .I(N__18961));
    LocalMux I__3255 (
            .O(N__18992),
            .I(N__18956));
    LocalMux I__3254 (
            .O(N__18989),
            .I(N__18956));
    Span4Mux_v I__3253 (
            .O(N__18980),
            .I(N__18953));
    LocalMux I__3252 (
            .O(N__18977),
            .I(N__18950));
    LocalMux I__3251 (
            .O(N__18972),
            .I(\processor_zipi8.t_state_1 ));
    Odrv4 I__3250 (
            .O(N__18969),
            .I(\processor_zipi8.t_state_1 ));
    LocalMux I__3249 (
            .O(N__18964),
            .I(\processor_zipi8.t_state_1 ));
    Odrv4 I__3248 (
            .O(N__18961),
            .I(\processor_zipi8.t_state_1 ));
    Odrv12 I__3247 (
            .O(N__18956),
            .I(\processor_zipi8.t_state_1 ));
    Odrv4 I__3246 (
            .O(N__18953),
            .I(\processor_zipi8.t_state_1 ));
    Odrv12 I__3245 (
            .O(N__18950),
            .I(\processor_zipi8.t_state_1 ));
    CascadeMux I__3244 (
            .O(N__18935),
            .I(\processor_zipi8.decode4_strobes_enables_i.register_enable_type_0_cascade_ ));
    CascadeMux I__3243 (
            .O(N__18932),
            .I(N__18922));
    CascadeMux I__3242 (
            .O(N__18931),
            .I(N__18918));
    CascadeMux I__3241 (
            .O(N__18930),
            .I(N__18915));
    CascadeMux I__3240 (
            .O(N__18929),
            .I(N__18909));
    InMux I__3239 (
            .O(N__18928),
            .I(N__18903));
    InMux I__3238 (
            .O(N__18927),
            .I(N__18903));
    InMux I__3237 (
            .O(N__18926),
            .I(N__18898));
    InMux I__3236 (
            .O(N__18925),
            .I(N__18898));
    InMux I__3235 (
            .O(N__18922),
            .I(N__18895));
    InMux I__3234 (
            .O(N__18921),
            .I(N__18890));
    InMux I__3233 (
            .O(N__18918),
            .I(N__18890));
    InMux I__3232 (
            .O(N__18915),
            .I(N__18885));
    InMux I__3231 (
            .O(N__18914),
            .I(N__18885));
    InMux I__3230 (
            .O(N__18913),
            .I(N__18880));
    InMux I__3229 (
            .O(N__18912),
            .I(N__18875));
    InMux I__3228 (
            .O(N__18909),
            .I(N__18875));
    CascadeMux I__3227 (
            .O(N__18908),
            .I(N__18871));
    LocalMux I__3226 (
            .O(N__18903),
            .I(N__18868));
    LocalMux I__3225 (
            .O(N__18898),
            .I(N__18863));
    LocalMux I__3224 (
            .O(N__18895),
            .I(N__18863));
    LocalMux I__3223 (
            .O(N__18890),
            .I(N__18858));
    LocalMux I__3222 (
            .O(N__18885),
            .I(N__18858));
    CascadeMux I__3221 (
            .O(N__18884),
            .I(N__18855));
    CascadeMux I__3220 (
            .O(N__18883),
            .I(N__18852));
    LocalMux I__3219 (
            .O(N__18880),
            .I(N__18849));
    LocalMux I__3218 (
            .O(N__18875),
            .I(N__18846));
    InMux I__3217 (
            .O(N__18874),
            .I(N__18841));
    InMux I__3216 (
            .O(N__18871),
            .I(N__18841));
    Span4Mux_v I__3215 (
            .O(N__18868),
            .I(N__18836));
    Span4Mux_v I__3214 (
            .O(N__18863),
            .I(N__18836));
    Span4Mux_s3_v I__3213 (
            .O(N__18858),
            .I(N__18833));
    InMux I__3212 (
            .O(N__18855),
            .I(N__18828));
    InMux I__3211 (
            .O(N__18852),
            .I(N__18828));
    Span4Mux_s2_h I__3210 (
            .O(N__18849),
            .I(N__18821));
    Span4Mux_h I__3209 (
            .O(N__18846),
            .I(N__18821));
    LocalMux I__3208 (
            .O(N__18841),
            .I(N__18821));
    Odrv4 I__3207 (
            .O(N__18836),
            .I(instruction_17));
    Odrv4 I__3206 (
            .O(N__18833),
            .I(instruction_17));
    LocalMux I__3205 (
            .O(N__18828),
            .I(instruction_17));
    Odrv4 I__3204 (
            .O(N__18821),
            .I(instruction_17));
    InMux I__3203 (
            .O(N__18812),
            .I(N__18806));
    InMux I__3202 (
            .O(N__18811),
            .I(N__18806));
    LocalMux I__3201 (
            .O(N__18806),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_22_3 ));
    InMux I__3200 (
            .O(N__18803),
            .I(N__18798));
    InMux I__3199 (
            .O(N__18802),
            .I(N__18794));
    InMux I__3198 (
            .O(N__18801),
            .I(N__18791));
    LocalMux I__3197 (
            .O(N__18798),
            .I(N__18788));
    InMux I__3196 (
            .O(N__18797),
            .I(N__18785));
    LocalMux I__3195 (
            .O(N__18794),
            .I(N__18778));
    LocalMux I__3194 (
            .O(N__18791),
            .I(N__18778));
    Span4Mux_v I__3193 (
            .O(N__18788),
            .I(N__18773));
    LocalMux I__3192 (
            .O(N__18785),
            .I(N__18773));
    CascadeMux I__3191 (
            .O(N__18784),
            .I(N__18770));
    CascadeMux I__3190 (
            .O(N__18783),
            .I(N__18767));
    Span4Mux_h I__3189 (
            .O(N__18778),
            .I(N__18762));
    Span4Mux_h I__3188 (
            .O(N__18773),
            .I(N__18759));
    InMux I__3187 (
            .O(N__18770),
            .I(N__18750));
    InMux I__3186 (
            .O(N__18767),
            .I(N__18750));
    InMux I__3185 (
            .O(N__18766),
            .I(N__18750));
    InMux I__3184 (
            .O(N__18765),
            .I(N__18750));
    Odrv4 I__3183 (
            .O(N__18762),
            .I(\processor_zipi8.sx_5 ));
    Odrv4 I__3182 (
            .O(N__18759),
            .I(\processor_zipi8.sx_5 ));
    LocalMux I__3181 (
            .O(N__18750),
            .I(\processor_zipi8.sx_5 ));
    InMux I__3180 (
            .O(N__18743),
            .I(N__18740));
    LocalMux I__3179 (
            .O(N__18740),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_4 ));
    CascadeMux I__3178 (
            .O(N__18737),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_4_cascade_ ));
    InMux I__3177 (
            .O(N__18734),
            .I(N__18731));
    LocalMux I__3176 (
            .O(N__18731),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_4 ));
    CascadeMux I__3175 (
            .O(N__18728),
            .I(N__18725));
    InMux I__3174 (
            .O(N__18725),
            .I(N__18719));
    InMux I__3173 (
            .O(N__18724),
            .I(N__18719));
    LocalMux I__3172 (
            .O(N__18719),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_4 ));
    InMux I__3171 (
            .O(N__18716),
            .I(N__18710));
    InMux I__3170 (
            .O(N__18715),
            .I(N__18710));
    LocalMux I__3169 (
            .O(N__18710),
            .I(N__18707));
    Span4Mux_h I__3168 (
            .O(N__18707),
            .I(N__18704));
    Odrv4 I__3167 (
            .O(N__18704),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_4 ));
    InMux I__3166 (
            .O(N__18701),
            .I(N__18695));
    InMux I__3165 (
            .O(N__18700),
            .I(N__18695));
    LocalMux I__3164 (
            .O(N__18695),
            .I(N__18692));
    Span4Mux_h I__3163 (
            .O(N__18692),
            .I(N__18689));
    Odrv4 I__3162 (
            .O(N__18689),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_4 ));
    CascadeMux I__3161 (
            .O(N__18686),
            .I(N__18682));
    InMux I__3160 (
            .O(N__18685),
            .I(N__18679));
    InMux I__3159 (
            .O(N__18682),
            .I(N__18676));
    LocalMux I__3158 (
            .O(N__18679),
            .I(N__18671));
    LocalMux I__3157 (
            .O(N__18676),
            .I(N__18671));
    Span12Mux_s9_v I__3156 (
            .O(N__18671),
            .I(N__18668));
    Odrv12 I__3155 (
            .O(N__18668),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_4 ));
    CascadeMux I__3154 (
            .O(N__18665),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_4_cascade_ ));
    InMux I__3153 (
            .O(N__18662),
            .I(N__18659));
    LocalMux I__3152 (
            .O(N__18659),
            .I(N__18656));
    Span4Mux_v I__3151 (
            .O(N__18656),
            .I(N__18653));
    Odrv4 I__3150 (
            .O(N__18653),
            .I(\processor_zipi8.shift_rotate_result_4 ));
    InMux I__3149 (
            .O(N__18650),
            .I(N__18647));
    LocalMux I__3148 (
            .O(N__18647),
            .I(N__18644));
    Span4Mux_h I__3147 (
            .O(N__18644),
            .I(N__18641));
    Odrv4 I__3146 (
            .O(N__18641),
            .I(\processor_zipi8.spm_data_4 ));
    CascadeMux I__3145 (
            .O(N__18638),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267_cascade_ ));
    InMux I__3144 (
            .O(N__18635),
            .I(N__18631));
    InMux I__3143 (
            .O(N__18634),
            .I(N__18628));
    LocalMux I__3142 (
            .O(N__18631),
            .I(N__18623));
    LocalMux I__3141 (
            .O(N__18628),
            .I(N__18623));
    Odrv4 I__3140 (
            .O(N__18623),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_4 ));
    CascadeMux I__3139 (
            .O(N__18620),
            .I(N__18617));
    InMux I__3138 (
            .O(N__18617),
            .I(N__18614));
    LocalMux I__3137 (
            .O(N__18614),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_4 ));
    InMux I__3136 (
            .O(N__18611),
            .I(N__18607));
    InMux I__3135 (
            .O(N__18610),
            .I(N__18604));
    LocalMux I__3134 (
            .O(N__18607),
            .I(N__18601));
    LocalMux I__3133 (
            .O(N__18604),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4 ));
    Odrv4 I__3132 (
            .O(N__18601),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4 ));
    InMux I__3131 (
            .O(N__18596),
            .I(N__18593));
    LocalMux I__3130 (
            .O(N__18593),
            .I(N__18590));
    Span4Mux_v I__3129 (
            .O(N__18590),
            .I(N__18587));
    Odrv4 I__3128 (
            .O(N__18587),
            .I(\processor_zipi8.shift_rotate_result_1 ));
    InMux I__3127 (
            .O(N__18584),
            .I(N__18581));
    LocalMux I__3126 (
            .O(N__18581),
            .I(N__18578));
    Span4Mux_h I__3125 (
            .O(N__18578),
            .I(N__18575));
    Odrv4 I__3124 (
            .O(N__18575),
            .I(\processor_zipi8.spm_data_1 ));
    CascadeMux I__3123 (
            .O(N__18572),
            .I(N__18568));
    InMux I__3122 (
            .O(N__18571),
            .I(N__18563));
    InMux I__3121 (
            .O(N__18568),
            .I(N__18563));
    LocalMux I__3120 (
            .O(N__18563),
            .I(N__18560));
    Odrv12 I__3119 (
            .O(N__18560),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_2 ));
    InMux I__3118 (
            .O(N__18557),
            .I(N__18553));
    InMux I__3117 (
            .O(N__18556),
            .I(N__18550));
    LocalMux I__3116 (
            .O(N__18553),
            .I(N__18545));
    LocalMux I__3115 (
            .O(N__18550),
            .I(N__18545));
    Span4Mux_v I__3114 (
            .O(N__18545),
            .I(N__18542));
    Odrv4 I__3113 (
            .O(N__18542),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_2 ));
    InMux I__3112 (
            .O(N__18539),
            .I(N__18536));
    LocalMux I__3111 (
            .O(N__18536),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_2 ));
    CascadeMux I__3110 (
            .O(N__18533),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_2_cascade_ ));
    CascadeMux I__3109 (
            .O(N__18530),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_2_cascade_ ));
    InMux I__3108 (
            .O(N__18527),
            .I(N__18524));
    LocalMux I__3107 (
            .O(N__18524),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_2 ));
    InMux I__3106 (
            .O(N__18521),
            .I(N__18517));
    InMux I__3105 (
            .O(N__18520),
            .I(N__18514));
    LocalMux I__3104 (
            .O(N__18517),
            .I(N__18511));
    LocalMux I__3103 (
            .O(N__18514),
            .I(N__18508));
    Span4Mux_v I__3102 (
            .O(N__18511),
            .I(N__18503));
    Span4Mux_v I__3101 (
            .O(N__18508),
            .I(N__18503));
    Span4Mux_h I__3100 (
            .O(N__18503),
            .I(N__18500));
    Odrv4 I__3099 (
            .O(N__18500),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_3 ));
    CascadeMux I__3098 (
            .O(N__18497),
            .I(N__18494));
    InMux I__3097 (
            .O(N__18494),
            .I(N__18491));
    LocalMux I__3096 (
            .O(N__18491),
            .I(N__18488));
    Odrv12 I__3095 (
            .O(N__18488),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_am_1_3 ));
    InMux I__3094 (
            .O(N__18485),
            .I(N__18481));
    InMux I__3093 (
            .O(N__18484),
            .I(N__18478));
    LocalMux I__3092 (
            .O(N__18481),
            .I(N__18475));
    LocalMux I__3091 (
            .O(N__18478),
            .I(N__18472));
    Span4Mux_h I__3090 (
            .O(N__18475),
            .I(N__18469));
    Span4Mux_h I__3089 (
            .O(N__18472),
            .I(N__18466));
    Odrv4 I__3088 (
            .O(N__18469),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3 ));
    Odrv4 I__3087 (
            .O(N__18466),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3 ));
    InMux I__3086 (
            .O(N__18461),
            .I(N__18458));
    LocalMux I__3085 (
            .O(N__18458),
            .I(N__18454));
    InMux I__3084 (
            .O(N__18457),
            .I(N__18451));
    Odrv4 I__3083 (
            .O(N__18454),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2 ));
    LocalMux I__3082 (
            .O(N__18451),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2 ));
    InMux I__3081 (
            .O(N__18446),
            .I(N__18442));
    InMux I__3080 (
            .O(N__18445),
            .I(N__18439));
    LocalMux I__3079 (
            .O(N__18442),
            .I(N__18436));
    LocalMux I__3078 (
            .O(N__18439),
            .I(N__18433));
    Span4Mux_h I__3077 (
            .O(N__18436),
            .I(N__18428));
    Span4Mux_v I__3076 (
            .O(N__18433),
            .I(N__18428));
    Odrv4 I__3075 (
            .O(N__18428),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_2 ));
    InMux I__3074 (
            .O(N__18425),
            .I(N__18422));
    LocalMux I__3073 (
            .O(N__18422),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_2 ));
    InMux I__3072 (
            .O(N__18419),
            .I(N__18413));
    InMux I__3071 (
            .O(N__18418),
            .I(N__18413));
    LocalMux I__3070 (
            .O(N__18413),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_4 ));
    CascadeMux I__3069 (
            .O(N__18410),
            .I(N__18406));
    InMux I__3068 (
            .O(N__18409),
            .I(N__18401));
    InMux I__3067 (
            .O(N__18406),
            .I(N__18401));
    LocalMux I__3066 (
            .O(N__18401),
            .I(N__18398));
    Span4Mux_v I__3065 (
            .O(N__18398),
            .I(N__18395));
    Odrv4 I__3064 (
            .O(N__18395),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_4 ));
    CascadeMux I__3063 (
            .O(N__18392),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_4_cascade_ ));
    CascadeMux I__3062 (
            .O(N__18389),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_2_cascade_ ));
    CascadeMux I__3061 (
            .O(N__18386),
            .I(N__18383));
    InMux I__3060 (
            .O(N__18383),
            .I(N__18379));
    InMux I__3059 (
            .O(N__18382),
            .I(N__18376));
    LocalMux I__3058 (
            .O(N__18379),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2 ));
    LocalMux I__3057 (
            .O(N__18376),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2 ));
    InMux I__3056 (
            .O(N__18371),
            .I(N__18365));
    InMux I__3055 (
            .O(N__18370),
            .I(N__18365));
    LocalMux I__3054 (
            .O(N__18365),
            .I(N__18362));
    Odrv4 I__3053 (
            .O(N__18362),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_2 ));
    InMux I__3052 (
            .O(N__18359),
            .I(N__18356));
    LocalMux I__3051 (
            .O(N__18356),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_bm_1_3 ));
    CascadeMux I__3050 (
            .O(N__18353),
            .I(N__18350));
    InMux I__3049 (
            .O(N__18350),
            .I(N__18344));
    InMux I__3048 (
            .O(N__18349),
            .I(N__18344));
    LocalMux I__3047 (
            .O(N__18344),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_3 ));
    InMux I__3046 (
            .O(N__18341),
            .I(N__18335));
    InMux I__3045 (
            .O(N__18340),
            .I(N__18335));
    LocalMux I__3044 (
            .O(N__18335),
            .I(N__18332));
    Odrv12 I__3043 (
            .O(N__18332),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_3 ));
    CascadeMux I__3042 (
            .O(N__18329),
            .I(N__18326));
    InMux I__3041 (
            .O(N__18326),
            .I(N__18322));
    InMux I__3040 (
            .O(N__18325),
            .I(N__18319));
    LocalMux I__3039 (
            .O(N__18322),
            .I(N__18314));
    LocalMux I__3038 (
            .O(N__18319),
            .I(N__18314));
    Span4Mux_h I__3037 (
            .O(N__18314),
            .I(N__18311));
    Odrv4 I__3036 (
            .O(N__18311),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_5 ));
    InMux I__3035 (
            .O(N__18308),
            .I(N__18302));
    InMux I__3034 (
            .O(N__18307),
            .I(N__18302));
    LocalMux I__3033 (
            .O(N__18302),
            .I(N__18299));
    Odrv4 I__3032 (
            .O(N__18299),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_5 ));
    InMux I__3031 (
            .O(N__18296),
            .I(N__18292));
    InMux I__3030 (
            .O(N__18295),
            .I(N__18289));
    LocalMux I__3029 (
            .O(N__18292),
            .I(N__18286));
    LocalMux I__3028 (
            .O(N__18289),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5 ));
    Odrv12 I__3027 (
            .O(N__18286),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5 ));
    CascadeMux I__3026 (
            .O(N__18281),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_5_cascade_ ));
    InMux I__3025 (
            .O(N__18278),
            .I(N__18275));
    LocalMux I__3024 (
            .O(N__18275),
            .I(N__18271));
    InMux I__3023 (
            .O(N__18274),
            .I(N__18268));
    Odrv12 I__3022 (
            .O(N__18271),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5 ));
    LocalMux I__3021 (
            .O(N__18268),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5 ));
    CascadeMux I__3020 (
            .O(N__18263),
            .I(N__18260));
    InMux I__3019 (
            .O(N__18260),
            .I(N__18257));
    LocalMux I__3018 (
            .O(N__18257),
            .I(N__18254));
    Span4Mux_v I__3017 (
            .O(N__18254),
            .I(N__18251));
    Span4Mux_h I__3016 (
            .O(N__18251),
            .I(N__18248));
    Odrv4 I__3015 (
            .O(N__18248),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_179 ));
    InMux I__3014 (
            .O(N__18245),
            .I(N__18239));
    InMux I__3013 (
            .O(N__18244),
            .I(N__18239));
    LocalMux I__3012 (
            .O(N__18239),
            .I(N__18236));
    Span4Mux_v I__3011 (
            .O(N__18236),
            .I(N__18233));
    Odrv4 I__3010 (
            .O(N__18233),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_2 ));
    CascadeMux I__3009 (
            .O(N__18230),
            .I(N__18227));
    InMux I__3008 (
            .O(N__18227),
            .I(N__18223));
    InMux I__3007 (
            .O(N__18226),
            .I(N__18220));
    LocalMux I__3006 (
            .O(N__18223),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2 ));
    LocalMux I__3005 (
            .O(N__18220),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2 ));
    CascadeMux I__3004 (
            .O(N__18215),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_2_cascade_ ));
    CascadeMux I__3003 (
            .O(N__18212),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_3_cascade_ ));
    InMux I__3002 (
            .O(N__18209),
            .I(N__18205));
    InMux I__3001 (
            .O(N__18208),
            .I(N__18202));
    LocalMux I__3000 (
            .O(N__18205),
            .I(N__18199));
    LocalMux I__2999 (
            .O(N__18202),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3 ));
    Odrv4 I__2998 (
            .O(N__18199),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3 ));
    InMux I__2997 (
            .O(N__18194),
            .I(N__18188));
    InMux I__2996 (
            .O(N__18193),
            .I(N__18188));
    LocalMux I__2995 (
            .O(N__18188),
            .I(N__18185));
    Odrv4 I__2994 (
            .O(N__18185),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_3 ));
    InMux I__2993 (
            .O(N__18182),
            .I(N__18179));
    LocalMux I__2992 (
            .O(N__18179),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_3 ));
    CascadeMux I__2991 (
            .O(N__18176),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_3_cascade_ ));
    InMux I__2990 (
            .O(N__18173),
            .I(N__18167));
    InMux I__2989 (
            .O(N__18172),
            .I(N__18167));
    LocalMux I__2988 (
            .O(N__18167),
            .I(N__18164));
    Odrv4 I__2987 (
            .O(N__18164),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_3 ));
    InMux I__2986 (
            .O(N__18161),
            .I(N__18155));
    InMux I__2985 (
            .O(N__18160),
            .I(N__18155));
    LocalMux I__2984 (
            .O(N__18155),
            .I(N__18152));
    Span4Mux_h I__2983 (
            .O(N__18152),
            .I(N__18149));
    Odrv4 I__2982 (
            .O(N__18149),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_3 ));
    InMux I__2981 (
            .O(N__18146),
            .I(N__18143));
    LocalMux I__2980 (
            .O(N__18143),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_3 ));
    InMux I__2979 (
            .O(N__18140),
            .I(N__18136));
    InMux I__2978 (
            .O(N__18139),
            .I(N__18133));
    LocalMux I__2977 (
            .O(N__18136),
            .I(N__18130));
    LocalMux I__2976 (
            .O(N__18133),
            .I(N__18127));
    Odrv4 I__2975 (
            .O(N__18130),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0 ));
    Odrv4 I__2974 (
            .O(N__18127),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0 ));
    CascadeMux I__2973 (
            .O(N__18122),
            .I(N__18118));
    CascadeMux I__2972 (
            .O(N__18121),
            .I(N__18115));
    InMux I__2971 (
            .O(N__18118),
            .I(N__18112));
    InMux I__2970 (
            .O(N__18115),
            .I(N__18109));
    LocalMux I__2969 (
            .O(N__18112),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0 ));
    LocalMux I__2968 (
            .O(N__18109),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0 ));
    InMux I__2967 (
            .O(N__18104),
            .I(N__18101));
    LocalMux I__2966 (
            .O(N__18101),
            .I(N__18098));
    Span4Mux_s2_h I__2965 (
            .O(N__18098),
            .I(N__18095));
    Span4Mux_h I__2964 (
            .O(N__18095),
            .I(N__18092));
    Odrv4 I__2963 (
            .O(N__18092),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_5 ));
    InMux I__2962 (
            .O(N__18089),
            .I(N__18086));
    LocalMux I__2961 (
            .O(N__18086),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_3 ));
    CEMux I__2960 (
            .O(N__18083),
            .I(N__18080));
    LocalMux I__2959 (
            .O(N__18080),
            .I(N__18077));
    Span4Mux_v I__2958 (
            .O(N__18077),
            .I(N__18073));
    CEMux I__2957 (
            .O(N__18076),
            .I(N__18070));
    Span4Mux_h I__2956 (
            .O(N__18073),
            .I(N__18067));
    LocalMux I__2955 (
            .O(N__18070),
            .I(N__18064));
    Sp12to4 I__2954 (
            .O(N__18067),
            .I(N__18059));
    Span12Mux_s3_v I__2953 (
            .O(N__18064),
            .I(N__18059));
    Odrv12 I__2952 (
            .O(N__18059),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe12 ));
    InMux I__2951 (
            .O(N__18056),
            .I(N__18053));
    LocalMux I__2950 (
            .O(N__18053),
            .I(\processor_zipi8.flags_i.use_zero_flagZ0 ));
    CascadeMux I__2949 (
            .O(N__18050),
            .I(\processor_zipi8.alu_result_0_cascade_ ));
    InMux I__2948 (
            .O(N__18047),
            .I(N__18044));
    LocalMux I__2947 (
            .O(N__18044),
            .I(N__18039));
    InMux I__2946 (
            .O(N__18043),
            .I(N__18034));
    InMux I__2945 (
            .O(N__18042),
            .I(N__18034));
    Span4Mux_v I__2944 (
            .O(N__18039),
            .I(N__18030));
    LocalMux I__2943 (
            .O(N__18034),
            .I(N__18026));
    InMux I__2942 (
            .O(N__18033),
            .I(N__18020));
    Span4Mux_v I__2941 (
            .O(N__18030),
            .I(N__18017));
    InMux I__2940 (
            .O(N__18029),
            .I(N__18014));
    Span4Mux_s2_v I__2939 (
            .O(N__18026),
            .I(N__18011));
    InMux I__2938 (
            .O(N__18025),
            .I(N__18004));
    InMux I__2937 (
            .O(N__18024),
            .I(N__18004));
    InMux I__2936 (
            .O(N__18023),
            .I(N__18004));
    LocalMux I__2935 (
            .O(N__18020),
            .I(\processor_zipi8.zero_flag ));
    Odrv4 I__2934 (
            .O(N__18017),
            .I(\processor_zipi8.zero_flag ));
    LocalMux I__2933 (
            .O(N__18014),
            .I(\processor_zipi8.zero_flag ));
    Odrv4 I__2932 (
            .O(N__18011),
            .I(\processor_zipi8.zero_flag ));
    LocalMux I__2931 (
            .O(N__18004),
            .I(\processor_zipi8.zero_flag ));
    CascadeMux I__2930 (
            .O(N__17993),
            .I(N__17985));
    InMux I__2929 (
            .O(N__17992),
            .I(N__17981));
    InMux I__2928 (
            .O(N__17991),
            .I(N__17978));
    InMux I__2927 (
            .O(N__17990),
            .I(N__17975));
    InMux I__2926 (
            .O(N__17989),
            .I(N__17971));
    InMux I__2925 (
            .O(N__17988),
            .I(N__17964));
    InMux I__2924 (
            .O(N__17985),
            .I(N__17964));
    InMux I__2923 (
            .O(N__17984),
            .I(N__17964));
    LocalMux I__2922 (
            .O(N__17981),
            .I(N__17961));
    LocalMux I__2921 (
            .O(N__17978),
            .I(N__17954));
    LocalMux I__2920 (
            .O(N__17975),
            .I(N__17954));
    InMux I__2919 (
            .O(N__17974),
            .I(N__17951));
    LocalMux I__2918 (
            .O(N__17971),
            .I(N__17946));
    LocalMux I__2917 (
            .O(N__17964),
            .I(N__17946));
    Span4Mux_h I__2916 (
            .O(N__17961),
            .I(N__17943));
    InMux I__2915 (
            .O(N__17960),
            .I(N__17938));
    InMux I__2914 (
            .O(N__17959),
            .I(N__17938));
    Span4Mux_v I__2913 (
            .O(N__17954),
            .I(N__17931));
    LocalMux I__2912 (
            .O(N__17951),
            .I(N__17931));
    Span4Mux_h I__2911 (
            .O(N__17946),
            .I(N__17931));
    Odrv4 I__2910 (
            .O(N__17943),
            .I(\processor_zipi8.carry_flag ));
    LocalMux I__2909 (
            .O(N__17938),
            .I(\processor_zipi8.carry_flag ));
    Odrv4 I__2908 (
            .O(N__17931),
            .I(\processor_zipi8.carry_flag ));
    InMux I__2907 (
            .O(N__17924),
            .I(N__17921));
    LocalMux I__2906 (
            .O(N__17921),
            .I(\processor_zipi8.N_11_0 ));
    InMux I__2905 (
            .O(N__17918),
            .I(N__17915));
    LocalMux I__2904 (
            .O(N__17915),
            .I(\processor_zipi8.alu_result_1 ));
    CascadeMux I__2903 (
            .O(N__17912),
            .I(\processor_zipi8.alu_result_2_cascade_ ));
    InMux I__2902 (
            .O(N__17909),
            .I(N__17906));
    LocalMux I__2901 (
            .O(N__17906),
            .I(\processor_zipi8.flags_i.zero_flag_3_0_0 ));
    InMux I__2900 (
            .O(N__17903),
            .I(N__17900));
    LocalMux I__2899 (
            .O(N__17900),
            .I(N__17897));
    Span4Mux_h I__2898 (
            .O(N__17897),
            .I(N__17894));
    Odrv4 I__2897 (
            .O(N__17894),
            .I(\processor_zipi8.flags_i.zero_flag_3_0_6 ));
    CascadeMux I__2896 (
            .O(N__17891),
            .I(N__17887));
    CascadeMux I__2895 (
            .O(N__17890),
            .I(N__17883));
    InMux I__2894 (
            .O(N__17887),
            .I(N__17872));
    InMux I__2893 (
            .O(N__17886),
            .I(N__17872));
    InMux I__2892 (
            .O(N__17883),
            .I(N__17872));
    InMux I__2891 (
            .O(N__17882),
            .I(N__17872));
    InMux I__2890 (
            .O(N__17881),
            .I(N__17868));
    LocalMux I__2889 (
            .O(N__17872),
            .I(N__17865));
    CascadeMux I__2888 (
            .O(N__17871),
            .I(N__17862));
    LocalMux I__2887 (
            .O(N__17868),
            .I(N__17854));
    Span4Mux_v I__2886 (
            .O(N__17865),
            .I(N__17851));
    InMux I__2885 (
            .O(N__17862),
            .I(N__17846));
    InMux I__2884 (
            .O(N__17861),
            .I(N__17841));
    InMux I__2883 (
            .O(N__17860),
            .I(N__17841));
    InMux I__2882 (
            .O(N__17859),
            .I(N__17834));
    InMux I__2881 (
            .O(N__17858),
            .I(N__17834));
    InMux I__2880 (
            .O(N__17857),
            .I(N__17834));
    Span4Mux_v I__2879 (
            .O(N__17854),
            .I(N__17831));
    Span4Mux_h I__2878 (
            .O(N__17851),
            .I(N__17828));
    InMux I__2877 (
            .O(N__17850),
            .I(N__17825));
    InMux I__2876 (
            .O(N__17849),
            .I(N__17822));
    LocalMux I__2875 (
            .O(N__17846),
            .I(N__17815));
    LocalMux I__2874 (
            .O(N__17841),
            .I(N__17815));
    LocalMux I__2873 (
            .O(N__17834),
            .I(N__17815));
    Odrv4 I__2872 (
            .O(N__17831),
            .I(\processor_zipi8.pc_mode_2 ));
    Odrv4 I__2871 (
            .O(N__17828),
            .I(\processor_zipi8.pc_mode_2 ));
    LocalMux I__2870 (
            .O(N__17825),
            .I(\processor_zipi8.pc_mode_2 ));
    LocalMux I__2869 (
            .O(N__17822),
            .I(\processor_zipi8.pc_mode_2 ));
    Odrv12 I__2868 (
            .O(N__17815),
            .I(\processor_zipi8.pc_mode_2 ));
    InMux I__2867 (
            .O(N__17804),
            .I(N__17795));
    InMux I__2866 (
            .O(N__17803),
            .I(N__17786));
    InMux I__2865 (
            .O(N__17802),
            .I(N__17786));
    InMux I__2864 (
            .O(N__17801),
            .I(N__17786));
    InMux I__2863 (
            .O(N__17800),
            .I(N__17786));
    InMux I__2862 (
            .O(N__17799),
            .I(N__17783));
    InMux I__2861 (
            .O(N__17798),
            .I(N__17780));
    LocalMux I__2860 (
            .O(N__17795),
            .I(N__17777));
    LocalMux I__2859 (
            .O(N__17786),
            .I(N__17768));
    LocalMux I__2858 (
            .O(N__17783),
            .I(N__17763));
    LocalMux I__2857 (
            .O(N__17780),
            .I(N__17763));
    Span4Mux_v I__2856 (
            .O(N__17777),
            .I(N__17760));
    InMux I__2855 (
            .O(N__17776),
            .I(N__17755));
    InMux I__2854 (
            .O(N__17775),
            .I(N__17755));
    InMux I__2853 (
            .O(N__17774),
            .I(N__17746));
    InMux I__2852 (
            .O(N__17773),
            .I(N__17746));
    InMux I__2851 (
            .O(N__17772),
            .I(N__17746));
    InMux I__2850 (
            .O(N__17771),
            .I(N__17746));
    Span4Mux_s1_h I__2849 (
            .O(N__17768),
            .I(N__17739));
    Span4Mux_h I__2848 (
            .O(N__17763),
            .I(N__17739));
    Span4Mux_h I__2847 (
            .O(N__17760),
            .I(N__17739));
    LocalMux I__2846 (
            .O(N__17755),
            .I(\processor_zipi8.pc_mode_1 ));
    LocalMux I__2845 (
            .O(N__17746),
            .I(\processor_zipi8.pc_mode_1 ));
    Odrv4 I__2844 (
            .O(N__17739),
            .I(\processor_zipi8.pc_mode_1 ));
    CascadeMux I__2843 (
            .O(N__17732),
            .I(N__17728));
    CascadeMux I__2842 (
            .O(N__17731),
            .I(N__17725));
    CascadeBuf I__2841 (
            .O(N__17728),
            .I(N__17722));
    CascadeBuf I__2840 (
            .O(N__17725),
            .I(N__17719));
    CascadeMux I__2839 (
            .O(N__17722),
            .I(N__17716));
    CascadeMux I__2838 (
            .O(N__17719),
            .I(N__17713));
    CascadeBuf I__2837 (
            .O(N__17716),
            .I(N__17710));
    CascadeBuf I__2836 (
            .O(N__17713),
            .I(N__17707));
    CascadeMux I__2835 (
            .O(N__17710),
            .I(N__17704));
    CascadeMux I__2834 (
            .O(N__17707),
            .I(N__17701));
    CascadeBuf I__2833 (
            .O(N__17704),
            .I(N__17698));
    CascadeBuf I__2832 (
            .O(N__17701),
            .I(N__17695));
    CascadeMux I__2831 (
            .O(N__17698),
            .I(N__17692));
    CascadeMux I__2830 (
            .O(N__17695),
            .I(N__17689));
    CascadeBuf I__2829 (
            .O(N__17692),
            .I(N__17686));
    CascadeBuf I__2828 (
            .O(N__17689),
            .I(N__17683));
    CascadeMux I__2827 (
            .O(N__17686),
            .I(N__17680));
    CascadeMux I__2826 (
            .O(N__17683),
            .I(N__17677));
    CascadeBuf I__2825 (
            .O(N__17680),
            .I(N__17674));
    CascadeBuf I__2824 (
            .O(N__17677),
            .I(N__17671));
    CascadeMux I__2823 (
            .O(N__17674),
            .I(N__17668));
    CascadeMux I__2822 (
            .O(N__17671),
            .I(N__17665));
    CascadeBuf I__2821 (
            .O(N__17668),
            .I(N__17662));
    CascadeBuf I__2820 (
            .O(N__17665),
            .I(N__17659));
    CascadeMux I__2819 (
            .O(N__17662),
            .I(N__17656));
    CascadeMux I__2818 (
            .O(N__17659),
            .I(N__17653));
    CascadeBuf I__2817 (
            .O(N__17656),
            .I(N__17650));
    CascadeBuf I__2816 (
            .O(N__17653),
            .I(N__17647));
    CascadeMux I__2815 (
            .O(N__17650),
            .I(N__17644));
    CascadeMux I__2814 (
            .O(N__17647),
            .I(N__17641));
    InMux I__2813 (
            .O(N__17644),
            .I(N__17636));
    InMux I__2812 (
            .O(N__17641),
            .I(N__17633));
    CascadeMux I__2811 (
            .O(N__17640),
            .I(N__17630));
    CascadeMux I__2810 (
            .O(N__17639),
            .I(N__17627));
    LocalMux I__2809 (
            .O(N__17636),
            .I(N__17624));
    LocalMux I__2808 (
            .O(N__17633),
            .I(N__17621));
    InMux I__2807 (
            .O(N__17630),
            .I(N__17617));
    InMux I__2806 (
            .O(N__17627),
            .I(N__17614));
    Span4Mux_s2_v I__2805 (
            .O(N__17624),
            .I(N__17609));
    Span4Mux_s2_v I__2804 (
            .O(N__17621),
            .I(N__17609));
    CascadeMux I__2803 (
            .O(N__17620),
            .I(N__17605));
    LocalMux I__2802 (
            .O(N__17617),
            .I(N__17602));
    LocalMux I__2801 (
            .O(N__17614),
            .I(N__17599));
    Span4Mux_h I__2800 (
            .O(N__17609),
            .I(N__17596));
    InMux I__2799 (
            .O(N__17608),
            .I(N__17593));
    InMux I__2798 (
            .O(N__17605),
            .I(N__17590));
    Span4Mux_v I__2797 (
            .O(N__17602),
            .I(N__17585));
    Span4Mux_h I__2796 (
            .O(N__17599),
            .I(N__17585));
    Span4Mux_v I__2795 (
            .O(N__17596),
            .I(N__17582));
    LocalMux I__2794 (
            .O(N__17593),
            .I(address_3));
    LocalMux I__2793 (
            .O(N__17590),
            .I(address_3));
    Odrv4 I__2792 (
            .O(N__17585),
            .I(address_3));
    Odrv4 I__2791 (
            .O(N__17582),
            .I(address_3));
    InMux I__2790 (
            .O(N__17573),
            .I(N__17570));
    LocalMux I__2789 (
            .O(N__17570),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_3 ));
    InMux I__2788 (
            .O(N__17567),
            .I(N__17564));
    LocalMux I__2787 (
            .O(N__17564),
            .I(N__17560));
    InMux I__2786 (
            .O(N__17563),
            .I(N__17557));
    Odrv4 I__2785 (
            .O(N__17560),
            .I(\processor_zipi8.arith_carry_in_0 ));
    LocalMux I__2784 (
            .O(N__17557),
            .I(\processor_zipi8.arith_carry_in_0 ));
    InMux I__2783 (
            .O(N__17552),
            .I(N__17549));
    LocalMux I__2782 (
            .O(N__17549),
            .I(N__17546));
    Odrv4 I__2781 (
            .O(N__17546),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0 ));
    InMux I__2780 (
            .O(N__17543),
            .I(N__17539));
    InMux I__2779 (
            .O(N__17542),
            .I(N__17536));
    LocalMux I__2778 (
            .O(N__17539),
            .I(N__17531));
    LocalMux I__2777 (
            .O(N__17536),
            .I(N__17531));
    Span4Mux_v I__2776 (
            .O(N__17531),
            .I(N__17527));
    InMux I__2775 (
            .O(N__17530),
            .I(N__17524));
    Odrv4 I__2774 (
            .O(N__17527),
            .I(\processor_zipi8.returni_type_o_2 ));
    LocalMux I__2773 (
            .O(N__17524),
            .I(\processor_zipi8.returni_type_o_2 ));
    InMux I__2772 (
            .O(N__17519),
            .I(N__17516));
    LocalMux I__2771 (
            .O(N__17516),
            .I(\processor_zipi8.decode4_strobes_enables_i.flag_enable_type_3 ));
    CascadeMux I__2770 (
            .O(N__17513),
            .I(\processor_zipi8.decode4_strobes_enables_i.un9_flag_enable_type_cascade_ ));
    CascadeMux I__2769 (
            .O(N__17510),
            .I(\processor_zipi8.decode4_strobes_enables_i.flag_enable_type_0_cascade_ ));
    CascadeMux I__2768 (
            .O(N__17507),
            .I(N__17503));
    InMux I__2767 (
            .O(N__17506),
            .I(N__17500));
    InMux I__2766 (
            .O(N__17503),
            .I(N__17497));
    LocalMux I__2765 (
            .O(N__17500),
            .I(N__17494));
    LocalMux I__2764 (
            .O(N__17497),
            .I(N__17491));
    Span4Mux_s1_h I__2763 (
            .O(N__17494),
            .I(N__17488));
    Odrv12 I__2762 (
            .O(N__17491),
            .I(\processor_zipi8.flag_enable ));
    Odrv4 I__2761 (
            .O(N__17488),
            .I(\processor_zipi8.flag_enable ));
    InMux I__2760 (
            .O(N__17483),
            .I(N__17480));
    LocalMux I__2759 (
            .O(N__17480),
            .I(\processor_zipi8.decode4_strobes_enables_i.spm_enable_value_1 ));
    CEMux I__2758 (
            .O(N__17477),
            .I(N__17474));
    LocalMux I__2757 (
            .O(N__17474),
            .I(N__17471));
    Span4Mux_v I__2756 (
            .O(N__17471),
            .I(N__17468));
    IoSpan4Mux I__2755 (
            .O(N__17468),
            .I(N__17465));
    IoSpan4Mux I__2754 (
            .O(N__17465),
            .I(N__17462));
    Span4Mux_s0_h I__2753 (
            .O(N__17462),
            .I(N__17459));
    Span4Mux_h I__2752 (
            .O(N__17459),
            .I(N__17456));
    Odrv4 I__2751 (
            .O(N__17456),
            .I(\processor_zipi8.spm_enable ));
    InMux I__2750 (
            .O(N__17453),
            .I(N__17450));
    LocalMux I__2749 (
            .O(N__17450),
            .I(N__17447));
    Odrv4 I__2748 (
            .O(N__17447),
            .I(\processor_zipi8.flags_i.carry_flag_value_1_0 ));
    SRMux I__2747 (
            .O(N__17444),
            .I(N__17438));
    InMux I__2746 (
            .O(N__17443),
            .I(N__17435));
    InMux I__2745 (
            .O(N__17442),
            .I(N__17430));
    InMux I__2744 (
            .O(N__17441),
            .I(N__17430));
    LocalMux I__2743 (
            .O(N__17438),
            .I(N__17426));
    LocalMux I__2742 (
            .O(N__17435),
            .I(N__17420));
    LocalMux I__2741 (
            .O(N__17430),
            .I(N__17420));
    SRMux I__2740 (
            .O(N__17429),
            .I(N__17417));
    Span4Mux_v I__2739 (
            .O(N__17426),
            .I(N__17409));
    SRMux I__2738 (
            .O(N__17425),
            .I(N__17406));
    Span4Mux_v I__2737 (
            .O(N__17420),
            .I(N__17395));
    LocalMux I__2736 (
            .O(N__17417),
            .I(N__17395));
    CascadeMux I__2735 (
            .O(N__17416),
            .I(N__17391));
    SRMux I__2734 (
            .O(N__17415),
            .I(N__17387));
    InMux I__2733 (
            .O(N__17414),
            .I(N__17380));
    InMux I__2732 (
            .O(N__17413),
            .I(N__17380));
    InMux I__2731 (
            .O(N__17412),
            .I(N__17380));
    Span4Mux_h I__2730 (
            .O(N__17409),
            .I(N__17374));
    LocalMux I__2729 (
            .O(N__17406),
            .I(N__17374));
    InMux I__2728 (
            .O(N__17405),
            .I(N__17365));
    InMux I__2727 (
            .O(N__17404),
            .I(N__17365));
    InMux I__2726 (
            .O(N__17403),
            .I(N__17365));
    InMux I__2725 (
            .O(N__17402),
            .I(N__17365));
    SRMux I__2724 (
            .O(N__17401),
            .I(N__17362));
    InMux I__2723 (
            .O(N__17400),
            .I(N__17359));
    Span4Mux_h I__2722 (
            .O(N__17395),
            .I(N__17356));
    InMux I__2721 (
            .O(N__17394),
            .I(N__17351));
    InMux I__2720 (
            .O(N__17391),
            .I(N__17351));
    SRMux I__2719 (
            .O(N__17390),
            .I(N__17348));
    LocalMux I__2718 (
            .O(N__17387),
            .I(N__17345));
    LocalMux I__2717 (
            .O(N__17380),
            .I(N__17342));
    CascadeMux I__2716 (
            .O(N__17379),
            .I(N__17336));
    Span4Mux_s2_h I__2715 (
            .O(N__17374),
            .I(N__17331));
    LocalMux I__2714 (
            .O(N__17365),
            .I(N__17331));
    LocalMux I__2713 (
            .O(N__17362),
            .I(N__17322));
    LocalMux I__2712 (
            .O(N__17359),
            .I(N__17322));
    Sp12to4 I__2711 (
            .O(N__17356),
            .I(N__17322));
    LocalMux I__2710 (
            .O(N__17351),
            .I(N__17322));
    LocalMux I__2709 (
            .O(N__17348),
            .I(N__17315));
    Span4Mux_v I__2708 (
            .O(N__17345),
            .I(N__17315));
    Span4Mux_v I__2707 (
            .O(N__17342),
            .I(N__17315));
    InMux I__2706 (
            .O(N__17341),
            .I(N__17308));
    InMux I__2705 (
            .O(N__17340),
            .I(N__17308));
    InMux I__2704 (
            .O(N__17339),
            .I(N__17308));
    InMux I__2703 (
            .O(N__17336),
            .I(N__17305));
    Span4Mux_s3_v I__2702 (
            .O(N__17331),
            .I(N__17302));
    Span12Mux_s6_v I__2701 (
            .O(N__17322),
            .I(N__17299));
    Span4Mux_h I__2700 (
            .O(N__17315),
            .I(N__17296));
    LocalMux I__2699 (
            .O(N__17308),
            .I(\processor_zipi8.internal_reset ));
    LocalMux I__2698 (
            .O(N__17305),
            .I(\processor_zipi8.internal_reset ));
    Odrv4 I__2697 (
            .O(N__17302),
            .I(\processor_zipi8.internal_reset ));
    Odrv12 I__2696 (
            .O(N__17299),
            .I(\processor_zipi8.internal_reset ));
    Odrv4 I__2695 (
            .O(N__17296),
            .I(\processor_zipi8.internal_reset ));
    InMux I__2694 (
            .O(N__17285),
            .I(N__17282));
    LocalMux I__2693 (
            .O(N__17282),
            .I(N__17278));
    InMux I__2692 (
            .O(N__17281),
            .I(N__17275));
    Span4Mux_h I__2691 (
            .O(N__17278),
            .I(N__17270));
    LocalMux I__2690 (
            .O(N__17275),
            .I(N__17270));
    Span4Mux_h I__2689 (
            .O(N__17270),
            .I(N__17267));
    Span4Mux_v I__2688 (
            .O(N__17267),
            .I(N__17264));
    Odrv4 I__2687 (
            .O(N__17264),
            .I(\processor_zipi8.flags_i.N_69 ));
    CascadeMux I__2686 (
            .O(N__17261),
            .I(N__17256));
    InMux I__2685 (
            .O(N__17260),
            .I(N__17252));
    CascadeMux I__2684 (
            .O(N__17259),
            .I(N__17248));
    InMux I__2683 (
            .O(N__17256),
            .I(N__17245));
    InMux I__2682 (
            .O(N__17255),
            .I(N__17242));
    LocalMux I__2681 (
            .O(N__17252),
            .I(N__17239));
    InMux I__2680 (
            .O(N__17251),
            .I(N__17234));
    InMux I__2679 (
            .O(N__17248),
            .I(N__17234));
    LocalMux I__2678 (
            .O(N__17245),
            .I(N__17231));
    LocalMux I__2677 (
            .O(N__17242),
            .I(N__17227));
    Sp12to4 I__2676 (
            .O(N__17239),
            .I(N__17222));
    LocalMux I__2675 (
            .O(N__17234),
            .I(N__17222));
    Span4Mux_v I__2674 (
            .O(N__17231),
            .I(N__17219));
    InMux I__2673 (
            .O(N__17230),
            .I(N__17216));
    Span12Mux_s11_v I__2672 (
            .O(N__17227),
            .I(N__17211));
    Span12Mux_s4_v I__2671 (
            .O(N__17222),
            .I(N__17211));
    Odrv4 I__2670 (
            .O(N__17219),
            .I(\processor_zipi8.stack_pointer_3 ));
    LocalMux I__2669 (
            .O(N__17216),
            .I(\processor_zipi8.stack_pointer_3 ));
    Odrv12 I__2668 (
            .O(N__17211),
            .I(\processor_zipi8.stack_pointer_3 ));
    CascadeMux I__2667 (
            .O(N__17204),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_3_cascade_ ));
    InMux I__2666 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__2665 (
            .O(N__17198),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_3 ));
    CascadeMux I__2664 (
            .O(N__17195),
            .I(\processor_zipi8.port_id_3_cascade_ ));
    InMux I__2663 (
            .O(N__17192),
            .I(N__17189));
    LocalMux I__2662 (
            .O(N__17189),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_3 ));
    CascadeMux I__2661 (
            .O(N__17186),
            .I(N__17182));
    CascadeMux I__2660 (
            .O(N__17185),
            .I(N__17179));
    InMux I__2659 (
            .O(N__17182),
            .I(N__17176));
    InMux I__2658 (
            .O(N__17179),
            .I(N__17173));
    LocalMux I__2657 (
            .O(N__17176),
            .I(N__17170));
    LocalMux I__2656 (
            .O(N__17173),
            .I(N__17167));
    Span4Mux_h I__2655 (
            .O(N__17170),
            .I(N__17163));
    Span4Mux_h I__2654 (
            .O(N__17167),
            .I(N__17160));
    CascadeMux I__2653 (
            .O(N__17166),
            .I(N__17157));
    Span4Mux_v I__2652 (
            .O(N__17163),
            .I(N__17152));
    Sp12to4 I__2651 (
            .O(N__17160),
            .I(N__17149));
    InMux I__2650 (
            .O(N__17157),
            .I(N__17142));
    InMux I__2649 (
            .O(N__17156),
            .I(N__17142));
    InMux I__2648 (
            .O(N__17155),
            .I(N__17142));
    Odrv4 I__2647 (
            .O(N__17152),
            .I(\processor_zipi8.port_id_3 ));
    Odrv12 I__2646 (
            .O(N__17149),
            .I(\processor_zipi8.port_id_3 ));
    LocalMux I__2645 (
            .O(N__17142),
            .I(\processor_zipi8.port_id_3 ));
    InMux I__2644 (
            .O(N__17135),
            .I(N__17132));
    LocalMux I__2643 (
            .O(N__17132),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_3 ));
    InMux I__2642 (
            .O(N__17129),
            .I(N__17110));
    InMux I__2641 (
            .O(N__17128),
            .I(N__17110));
    InMux I__2640 (
            .O(N__17127),
            .I(N__17110));
    InMux I__2639 (
            .O(N__17126),
            .I(N__17110));
    InMux I__2638 (
            .O(N__17125),
            .I(N__17110));
    InMux I__2637 (
            .O(N__17124),
            .I(N__17103));
    InMux I__2636 (
            .O(N__17123),
            .I(N__17103));
    InMux I__2635 (
            .O(N__17122),
            .I(N__17103));
    InMux I__2634 (
            .O(N__17121),
            .I(N__17097));
    LocalMux I__2633 (
            .O(N__17110),
            .I(N__17092));
    LocalMux I__2632 (
            .O(N__17103),
            .I(N__17092));
    InMux I__2631 (
            .O(N__17102),
            .I(N__17089));
    InMux I__2630 (
            .O(N__17101),
            .I(N__17084));
    InMux I__2629 (
            .O(N__17100),
            .I(N__17084));
    LocalMux I__2628 (
            .O(N__17097),
            .I(N__17077));
    Span4Mux_h I__2627 (
            .O(N__17092),
            .I(N__17077));
    LocalMux I__2626 (
            .O(N__17089),
            .I(N__17077));
    LocalMux I__2625 (
            .O(N__17084),
            .I(N__17074));
    Span4Mux_v I__2624 (
            .O(N__17077),
            .I(N__17071));
    Span4Mux_h I__2623 (
            .O(N__17074),
            .I(N__17068));
    Sp12to4 I__2622 (
            .O(N__17071),
            .I(N__17065));
    Sp12to4 I__2621 (
            .O(N__17068),
            .I(N__17062));
    Span12Mux_s2_h I__2620 (
            .O(N__17065),
            .I(N__17057));
    Span12Mux_v I__2619 (
            .O(N__17062),
            .I(N__17057));
    Odrv12 I__2618 (
            .O(N__17057),
            .I(instruction_3));
    InMux I__2617 (
            .O(N__17054),
            .I(N__17051));
    LocalMux I__2616 (
            .O(N__17051),
            .I(\processor_zipi8.pc_vector_3 ));
    CascadeMux I__2615 (
            .O(N__17048),
            .I(N__17045));
    InMux I__2614 (
            .O(N__17045),
            .I(N__17042));
    LocalMux I__2613 (
            .O(N__17042),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_0 ));
    InMux I__2612 (
            .O(N__17039),
            .I(N__17036));
    LocalMux I__2611 (
            .O(N__17036),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4Z0Z_0 ));
    CascadeMux I__2610 (
            .O(N__17033),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_cascade_ ));
    InMux I__2609 (
            .O(N__17030),
            .I(N__17027));
    LocalMux I__2608 (
            .O(N__17027),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0 ));
    CascadeMux I__2607 (
            .O(N__17024),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0_cascade_ ));
    InMux I__2606 (
            .O(N__17021),
            .I(N__17018));
    LocalMux I__2605 (
            .O(N__17018),
            .I(N__17015));
    Span4Mux_h I__2604 (
            .O(N__17015),
            .I(N__17011));
    InMux I__2603 (
            .O(N__17014),
            .I(N__17008));
    Odrv4 I__2602 (
            .O(N__17011),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1 ));
    LocalMux I__2601 (
            .O(N__17008),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1 ));
    InMux I__2600 (
            .O(N__17003),
            .I(N__16997));
    InMux I__2599 (
            .O(N__17002),
            .I(N__16994));
    InMux I__2598 (
            .O(N__17001),
            .I(N__16989));
    InMux I__2597 (
            .O(N__17000),
            .I(N__16989));
    LocalMux I__2596 (
            .O(N__16997),
            .I(N__16984));
    LocalMux I__2595 (
            .O(N__16994),
            .I(N__16984));
    LocalMux I__2594 (
            .O(N__16989),
            .I(N__16981));
    Span4Mux_v I__2593 (
            .O(N__16984),
            .I(N__16976));
    Span4Mux_v I__2592 (
            .O(N__16981),
            .I(N__16976));
    Span4Mux_h I__2591 (
            .O(N__16976),
            .I(N__16973));
    Span4Mux_v I__2590 (
            .O(N__16973),
            .I(N__16970));
    Span4Mux_v I__2589 (
            .O(N__16970),
            .I(N__16967));
    Odrv4 I__2588 (
            .O(N__16967),
            .I(instruction_0));
    InMux I__2587 (
            .O(N__16964),
            .I(N__16961));
    LocalMux I__2586 (
            .O(N__16961),
            .I(N__16958));
    Span4Mux_h I__2585 (
            .O(N__16958),
            .I(N__16955));
    Odrv4 I__2584 (
            .O(N__16955),
            .I(\processor_zipi8.register_bank_control_i.un1_bank_value ));
    CascadeMux I__2583 (
            .O(N__16952),
            .I(\processor_zipi8.register_bank_control_i.bank_0_1_cascade_ ));
    InMux I__2582 (
            .O(N__16949),
            .I(N__16945));
    InMux I__2581 (
            .O(N__16948),
            .I(N__16942));
    LocalMux I__2580 (
            .O(N__16945),
            .I(N__16939));
    LocalMux I__2579 (
            .O(N__16942),
            .I(N__16936));
    Odrv12 I__2578 (
            .O(N__16939),
            .I(\processor_zipi8.sy_4 ));
    Odrv4 I__2577 (
            .O(N__16936),
            .I(\processor_zipi8.sy_4 ));
    InMux I__2576 (
            .O(N__16931),
            .I(N__16928));
    LocalMux I__2575 (
            .O(N__16928),
            .I(N__16925));
    Span4Mux_h I__2574 (
            .O(N__16925),
            .I(N__16922));
    Span4Mux_s2_h I__2573 (
            .O(N__16922),
            .I(N__16919));
    Odrv4 I__2572 (
            .O(N__16919),
            .I(\processor_zipi8.stack_i.stack_bank ));
    InMux I__2571 (
            .O(N__16916),
            .I(N__16913));
    LocalMux I__2570 (
            .O(N__16913),
            .I(\processor_zipi8.shadow_bank ));
    InMux I__2569 (
            .O(N__16910),
            .I(N__16907));
    LocalMux I__2568 (
            .O(N__16907),
            .I(N__16904));
    Span4Mux_h I__2567 (
            .O(N__16904),
            .I(N__16900));
    InMux I__2566 (
            .O(N__16903),
            .I(N__16897));
    Odrv4 I__2565 (
            .O(N__16900),
            .I(\processor_zipi8.un16_alu_mux_sel_value ));
    LocalMux I__2564 (
            .O(N__16897),
            .I(\processor_zipi8.un16_alu_mux_sel_value ));
    CascadeMux I__2563 (
            .O(N__16892),
            .I(\processor_zipi8.un4_arith_logical_sel_cascade_ ));
    InMux I__2562 (
            .O(N__16889),
            .I(N__16886));
    LocalMux I__2561 (
            .O(N__16886),
            .I(N__16883));
    Span4Mux_s2_h I__2560 (
            .O(N__16883),
            .I(N__16880));
    Span4Mux_v I__2559 (
            .O(N__16880),
            .I(N__16876));
    InMux I__2558 (
            .O(N__16879),
            .I(N__16873));
    Odrv4 I__2557 (
            .O(N__16876),
            .I(\processor_zipi8.alu_mux_sel_value_1 ));
    LocalMux I__2556 (
            .O(N__16873),
            .I(\processor_zipi8.alu_mux_sel_value_1 ));
    InMux I__2555 (
            .O(N__16868),
            .I(N__16865));
    LocalMux I__2554 (
            .O(N__16865),
            .I(N__16862));
    Span4Mux_v I__2553 (
            .O(N__16862),
            .I(N__16858));
    InMux I__2552 (
            .O(N__16861),
            .I(N__16855));
    Odrv4 I__2551 (
            .O(N__16858),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2 ));
    LocalMux I__2550 (
            .O(N__16855),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2 ));
    CascadeMux I__2549 (
            .O(N__16850),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2_cascade_ ));
    CascadeMux I__2548 (
            .O(N__16847),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_0_cascade_ ));
    CascadeMux I__2547 (
            .O(N__16844),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_0_cascade_ ));
    CascadeMux I__2546 (
            .O(N__16841),
            .I(N__16837));
    CascadeMux I__2545 (
            .O(N__16840),
            .I(N__16834));
    InMux I__2544 (
            .O(N__16837),
            .I(N__16831));
    InMux I__2543 (
            .O(N__16834),
            .I(N__16828));
    LocalMux I__2542 (
            .O(N__16831),
            .I(N__16825));
    LocalMux I__2541 (
            .O(N__16828),
            .I(N__16816));
    Span4Mux_s3_h I__2540 (
            .O(N__16825),
            .I(N__16816));
    InMux I__2539 (
            .O(N__16824),
            .I(N__16811));
    InMux I__2538 (
            .O(N__16823),
            .I(N__16811));
    InMux I__2537 (
            .O(N__16822),
            .I(N__16806));
    InMux I__2536 (
            .O(N__16821),
            .I(N__16806));
    Odrv4 I__2535 (
            .O(N__16816),
            .I(\processor_zipi8.port_id_0 ));
    LocalMux I__2534 (
            .O(N__16811),
            .I(\processor_zipi8.port_id_0 ));
    LocalMux I__2533 (
            .O(N__16806),
            .I(\processor_zipi8.port_id_0 ));
    InMux I__2532 (
            .O(N__16799),
            .I(N__16793));
    InMux I__2531 (
            .O(N__16798),
            .I(N__16793));
    LocalMux I__2530 (
            .O(N__16793),
            .I(N__16790));
    Span4Mux_h I__2529 (
            .O(N__16790),
            .I(N__16787));
    Odrv4 I__2528 (
            .O(N__16787),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_6 ));
    CascadeMux I__2527 (
            .O(N__16784),
            .I(\processor_zipi8.flags_i.carry_flag_value_1_1_cascade_ ));
    InMux I__2526 (
            .O(N__16781),
            .I(N__16778));
    LocalMux I__2525 (
            .O(N__16778),
            .I(\processor_zipi8.flags_i.parity_4 ));
    InMux I__2524 (
            .O(N__16775),
            .I(N__16772));
    LocalMux I__2523 (
            .O(N__16772),
            .I(\processor_zipi8.flags_i.carry_flag_RNOZ0Z_1 ));
    InMux I__2522 (
            .O(N__16769),
            .I(N__16765));
    InMux I__2521 (
            .O(N__16768),
            .I(N__16762));
    LocalMux I__2520 (
            .O(N__16765),
            .I(\processor_zipi8.flags_i.arith_carryZ0 ));
    LocalMux I__2519 (
            .O(N__16762),
            .I(\processor_zipi8.flags_i.arith_carryZ0 ));
    CascadeMux I__2518 (
            .O(N__16757),
            .I(N__16753));
    InMux I__2517 (
            .O(N__16756),
            .I(N__16748));
    InMux I__2516 (
            .O(N__16753),
            .I(N__16748));
    LocalMux I__2515 (
            .O(N__16748),
            .I(N__16745));
    Span4Mux_v I__2514 (
            .O(N__16745),
            .I(N__16742));
    Span4Mux_h I__2513 (
            .O(N__16742),
            .I(N__16739));
    Odrv4 I__2512 (
            .O(N__16739),
            .I(\processor_zipi8.flags_i.shift_carryZ0 ));
    InMux I__2511 (
            .O(N__16736),
            .I(N__16733));
    LocalMux I__2510 (
            .O(N__16733),
            .I(\processor_zipi8.flags_i.carry_flag_value_1_0_0 ));
    InMux I__2509 (
            .O(N__16730),
            .I(N__16727));
    LocalMux I__2508 (
            .O(N__16727),
            .I(N__16724));
    Span4Mux_v I__2507 (
            .O(N__16724),
            .I(N__16721));
    Odrv4 I__2506 (
            .O(N__16721),
            .I(\processor_zipi8.decode4_pc_statck_i.N_22_0 ));
    InMux I__2505 (
            .O(N__16718),
            .I(N__16715));
    LocalMux I__2504 (
            .O(N__16715),
            .I(\processor_zipi8.register_bank_control_i.un17_regbank_type_1 ));
    InMux I__2503 (
            .O(N__16712),
            .I(N__16709));
    LocalMux I__2502 (
            .O(N__16709),
            .I(\processor_zipi8.flags_i.un17_carry_flag_value_0 ));
    CascadeMux I__2501 (
            .O(N__16706),
            .I(N__16703));
    InMux I__2500 (
            .O(N__16703),
            .I(N__16698));
    InMux I__2499 (
            .O(N__16702),
            .I(N__16695));
    InMux I__2498 (
            .O(N__16701),
            .I(N__16691));
    LocalMux I__2497 (
            .O(N__16698),
            .I(N__16686));
    LocalMux I__2496 (
            .O(N__16695),
            .I(N__16686));
    InMux I__2495 (
            .O(N__16694),
            .I(N__16680));
    LocalMux I__2494 (
            .O(N__16691),
            .I(N__16674));
    Span4Mux_v I__2493 (
            .O(N__16686),
            .I(N__16674));
    CascadeMux I__2492 (
            .O(N__16685),
            .I(N__16671));
    CascadeMux I__2491 (
            .O(N__16684),
            .I(N__16668));
    CascadeMux I__2490 (
            .O(N__16683),
            .I(N__16664));
    LocalMux I__2489 (
            .O(N__16680),
            .I(N__16661));
    InMux I__2488 (
            .O(N__16679),
            .I(N__16658));
    Span4Mux_h I__2487 (
            .O(N__16674),
            .I(N__16655));
    InMux I__2486 (
            .O(N__16671),
            .I(N__16648));
    InMux I__2485 (
            .O(N__16668),
            .I(N__16648));
    InMux I__2484 (
            .O(N__16667),
            .I(N__16648));
    InMux I__2483 (
            .O(N__16664),
            .I(N__16645));
    Odrv12 I__2482 (
            .O(N__16661),
            .I(\processor_zipi8.sx_7 ));
    LocalMux I__2481 (
            .O(N__16658),
            .I(\processor_zipi8.sx_7 ));
    Odrv4 I__2480 (
            .O(N__16655),
            .I(\processor_zipi8.sx_7 ));
    LocalMux I__2479 (
            .O(N__16648),
            .I(\processor_zipi8.sx_7 ));
    LocalMux I__2478 (
            .O(N__16645),
            .I(\processor_zipi8.sx_7 ));
    CascadeMux I__2477 (
            .O(N__16634),
            .I(N__16627));
    CascadeMux I__2476 (
            .O(N__16633),
            .I(N__16624));
    InMux I__2475 (
            .O(N__16632),
            .I(N__16620));
    CascadeMux I__2474 (
            .O(N__16631),
            .I(N__16616));
    InMux I__2473 (
            .O(N__16630),
            .I(N__16610));
    InMux I__2472 (
            .O(N__16627),
            .I(N__16610));
    InMux I__2471 (
            .O(N__16624),
            .I(N__16605));
    InMux I__2470 (
            .O(N__16623),
            .I(N__16605));
    LocalMux I__2469 (
            .O(N__16620),
            .I(N__16602));
    CascadeMux I__2468 (
            .O(N__16619),
            .I(N__16599));
    InMux I__2467 (
            .O(N__16616),
            .I(N__16594));
    InMux I__2466 (
            .O(N__16615),
            .I(N__16594));
    LocalMux I__2465 (
            .O(N__16610),
            .I(N__16589));
    LocalMux I__2464 (
            .O(N__16605),
            .I(N__16589));
    Span4Mux_v I__2463 (
            .O(N__16602),
            .I(N__16586));
    InMux I__2462 (
            .O(N__16599),
            .I(N__16583));
    LocalMux I__2461 (
            .O(N__16594),
            .I(N__16578));
    Span4Mux_h I__2460 (
            .O(N__16589),
            .I(N__16578));
    Span4Mux_s2_h I__2459 (
            .O(N__16586),
            .I(N__16575));
    LocalMux I__2458 (
            .O(N__16583),
            .I(N__16572));
    Span4Mux_v I__2457 (
            .O(N__16578),
            .I(N__16569));
    Odrv4 I__2456 (
            .O(N__16575),
            .I(\processor_zipi8.sx_6 ));
    Odrv12 I__2455 (
            .O(N__16572),
            .I(\processor_zipi8.sx_6 ));
    Odrv4 I__2454 (
            .O(N__16569),
            .I(\processor_zipi8.sx_6 ));
    InMux I__2453 (
            .O(N__16562),
            .I(N__16559));
    LocalMux I__2452 (
            .O(N__16559),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6 ));
    CascadeMux I__2451 (
            .O(N__16556),
            .I(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6_cascade_ ));
    InMux I__2450 (
            .O(N__16553),
            .I(N__16547));
    InMux I__2449 (
            .O(N__16552),
            .I(N__16547));
    LocalMux I__2448 (
            .O(N__16547),
            .I(N__16544));
    Odrv12 I__2447 (
            .O(N__16544),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_7 ));
    InMux I__2446 (
            .O(N__16541),
            .I(N__16538));
    LocalMux I__2445 (
            .O(N__16538),
            .I(N__16534));
    InMux I__2444 (
            .O(N__16537),
            .I(N__16531));
    Span4Mux_v I__2443 (
            .O(N__16534),
            .I(N__16526));
    LocalMux I__2442 (
            .O(N__16531),
            .I(N__16526));
    Odrv4 I__2441 (
            .O(N__16526),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_7 ));
    CEMux I__2440 (
            .O(N__16523),
            .I(N__16520));
    LocalMux I__2439 (
            .O(N__16520),
            .I(N__16517));
    Span4Mux_v I__2438 (
            .O(N__16517),
            .I(N__16514));
    Odrv4 I__2437 (
            .O(N__16514),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe15 ));
    CascadeMux I__2436 (
            .O(N__16511),
            .I(N__16507));
    InMux I__2435 (
            .O(N__16510),
            .I(N__16502));
    InMux I__2434 (
            .O(N__16507),
            .I(N__16502));
    LocalMux I__2433 (
            .O(N__16502),
            .I(N__16499));
    Odrv4 I__2432 (
            .O(N__16499),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_0 ));
    InMux I__2431 (
            .O(N__16496),
            .I(N__16490));
    InMux I__2430 (
            .O(N__16495),
            .I(N__16490));
    LocalMux I__2429 (
            .O(N__16490),
            .I(N__16487));
    Odrv12 I__2428 (
            .O(N__16487),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_5 ));
    InMux I__2427 (
            .O(N__16484),
            .I(N__16478));
    InMux I__2426 (
            .O(N__16483),
            .I(N__16478));
    LocalMux I__2425 (
            .O(N__16478),
            .I(N__16475));
    Span4Mux_h I__2424 (
            .O(N__16475),
            .I(N__16472));
    Odrv4 I__2423 (
            .O(N__16472),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_6 ));
    InMux I__2422 (
            .O(N__16469),
            .I(N__16463));
    InMux I__2421 (
            .O(N__16468),
            .I(N__16463));
    LocalMux I__2420 (
            .O(N__16463),
            .I(N__16460));
    Span4Mux_v I__2419 (
            .O(N__16460),
            .I(N__16457));
    Odrv4 I__2418 (
            .O(N__16457),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_7 ));
    CEMux I__2417 (
            .O(N__16454),
            .I(N__16451));
    LocalMux I__2416 (
            .O(N__16451),
            .I(N__16448));
    Odrv4 I__2415 (
            .O(N__16448),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe9 ));
    CascadeMux I__2414 (
            .O(N__16445),
            .I(N__16442));
    InMux I__2413 (
            .O(N__16442),
            .I(N__16436));
    InMux I__2412 (
            .O(N__16441),
            .I(N__16436));
    LocalMux I__2411 (
            .O(N__16436),
            .I(N__16433));
    Span4Mux_v I__2410 (
            .O(N__16433),
            .I(N__16430));
    Odrv4 I__2409 (
            .O(N__16430),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_6 ));
    InMux I__2408 (
            .O(N__16427),
            .I(N__16423));
    InMux I__2407 (
            .O(N__16426),
            .I(N__16420));
    LocalMux I__2406 (
            .O(N__16423),
            .I(N__16415));
    LocalMux I__2405 (
            .O(N__16420),
            .I(N__16415));
    Span4Mux_h I__2404 (
            .O(N__16415),
            .I(N__16412));
    Odrv4 I__2403 (
            .O(N__16412),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_7 ));
    CEMux I__2402 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__2401 (
            .O(N__16406),
            .I(N__16403));
    Span4Mux_v I__2400 (
            .O(N__16403),
            .I(N__16400));
    Span4Mux_s1_v I__2399 (
            .O(N__16400),
            .I(N__16397));
    Odrv4 I__2398 (
            .O(N__16397),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe13 ));
    InMux I__2397 (
            .O(N__16394),
            .I(N__16388));
    InMux I__2396 (
            .O(N__16393),
            .I(N__16388));
    LocalMux I__2395 (
            .O(N__16388),
            .I(N__16385));
    Span4Mux_v I__2394 (
            .O(N__16385),
            .I(N__16382));
    Odrv4 I__2393 (
            .O(N__16382),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_6 ));
    InMux I__2392 (
            .O(N__16379),
            .I(N__16375));
    InMux I__2391 (
            .O(N__16378),
            .I(N__16372));
    LocalMux I__2390 (
            .O(N__16375),
            .I(N__16369));
    LocalMux I__2389 (
            .O(N__16372),
            .I(N__16366));
    Odrv4 I__2388 (
            .O(N__16369),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6 ));
    Odrv12 I__2387 (
            .O(N__16366),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6 ));
    InMux I__2386 (
            .O(N__16361),
            .I(N__16357));
    InMux I__2385 (
            .O(N__16360),
            .I(N__16354));
    LocalMux I__2384 (
            .O(N__16357),
            .I(N__16349));
    LocalMux I__2383 (
            .O(N__16354),
            .I(N__16349));
    Odrv4 I__2382 (
            .O(N__16349),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_6 ));
    CascadeMux I__2381 (
            .O(N__16346),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_6_cascade_ ));
    InMux I__2380 (
            .O(N__16343),
            .I(N__16340));
    LocalMux I__2379 (
            .O(N__16340),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIK4HN1_6 ));
    InMux I__2378 (
            .O(N__16337),
            .I(N__16334));
    LocalMux I__2377 (
            .O(N__16334),
            .I(N__16331));
    Odrv4 I__2376 (
            .O(N__16331),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNII1NP1_6 ));
    InMux I__2375 (
            .O(N__16328),
            .I(N__16325));
    LocalMux I__2374 (
            .O(N__16325),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_6 ));
    CascadeMux I__2373 (
            .O(N__16322),
            .I(N__16319));
    InMux I__2372 (
            .O(N__16319),
            .I(N__16316));
    LocalMux I__2371 (
            .O(N__16316),
            .I(N__16313));
    Span4Mux_h I__2370 (
            .O(N__16313),
            .I(N__16310));
    Odrv4 I__2369 (
            .O(N__16310),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIGUSR1_6 ));
    CascadeMux I__2368 (
            .O(N__16307),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7B4G8_6_cascade_ ));
    InMux I__2367 (
            .O(N__16304),
            .I(N__16301));
    LocalMux I__2366 (
            .O(N__16301),
            .I(\processor_zipi8.decode4_pc_statck_i.un3_pc_modeZ0 ));
    InMux I__2365 (
            .O(N__16298),
            .I(N__16295));
    LocalMux I__2364 (
            .O(N__16295),
            .I(\processor_zipi8.N_17_0 ));
    CascadeMux I__2363 (
            .O(N__16292),
            .I(N__16284));
    CascadeMux I__2362 (
            .O(N__16291),
            .I(N__16281));
    CascadeMux I__2361 (
            .O(N__16290),
            .I(N__16272));
    InMux I__2360 (
            .O(N__16289),
            .I(N__16265));
    InMux I__2359 (
            .O(N__16288),
            .I(N__16265));
    InMux I__2358 (
            .O(N__16287),
            .I(N__16262));
    InMux I__2357 (
            .O(N__16284),
            .I(N__16259));
    InMux I__2356 (
            .O(N__16281),
            .I(N__16256));
    InMux I__2355 (
            .O(N__16280),
            .I(N__16253));
    InMux I__2354 (
            .O(N__16279),
            .I(N__16246));
    InMux I__2353 (
            .O(N__16278),
            .I(N__16246));
    InMux I__2352 (
            .O(N__16277),
            .I(N__16246));
    InMux I__2351 (
            .O(N__16276),
            .I(N__16237));
    InMux I__2350 (
            .O(N__16275),
            .I(N__16237));
    InMux I__2349 (
            .O(N__16272),
            .I(N__16237));
    InMux I__2348 (
            .O(N__16271),
            .I(N__16237));
    InMux I__2347 (
            .O(N__16270),
            .I(N__16234));
    LocalMux I__2346 (
            .O(N__16265),
            .I(N__16213));
    LocalMux I__2345 (
            .O(N__16262),
            .I(N__16210));
    LocalMux I__2344 (
            .O(N__16259),
            .I(N__16207));
    LocalMux I__2343 (
            .O(N__16256),
            .I(N__16204));
    LocalMux I__2342 (
            .O(N__16253),
            .I(N__16201));
    LocalMux I__2341 (
            .O(N__16246),
            .I(N__16198));
    LocalMux I__2340 (
            .O(N__16237),
            .I(N__16195));
    LocalMux I__2339 (
            .O(N__16234),
            .I(N__16192));
    CEMux I__2338 (
            .O(N__16233),
            .I(N__16139));
    CEMux I__2337 (
            .O(N__16232),
            .I(N__16139));
    CEMux I__2336 (
            .O(N__16231),
            .I(N__16139));
    CEMux I__2335 (
            .O(N__16230),
            .I(N__16139));
    CEMux I__2334 (
            .O(N__16229),
            .I(N__16139));
    CEMux I__2333 (
            .O(N__16228),
            .I(N__16139));
    CEMux I__2332 (
            .O(N__16227),
            .I(N__16139));
    CEMux I__2331 (
            .O(N__16226),
            .I(N__16139));
    CEMux I__2330 (
            .O(N__16225),
            .I(N__16139));
    CEMux I__2329 (
            .O(N__16224),
            .I(N__16139));
    CEMux I__2328 (
            .O(N__16223),
            .I(N__16139));
    CEMux I__2327 (
            .O(N__16222),
            .I(N__16139));
    CEMux I__2326 (
            .O(N__16221),
            .I(N__16139));
    CEMux I__2325 (
            .O(N__16220),
            .I(N__16139));
    CEMux I__2324 (
            .O(N__16219),
            .I(N__16139));
    CEMux I__2323 (
            .O(N__16218),
            .I(N__16139));
    CEMux I__2322 (
            .O(N__16217),
            .I(N__16139));
    CEMux I__2321 (
            .O(N__16216),
            .I(N__16139));
    Glb2LocalMux I__2320 (
            .O(N__16213),
            .I(N__16139));
    Glb2LocalMux I__2319 (
            .O(N__16210),
            .I(N__16139));
    Glb2LocalMux I__2318 (
            .O(N__16207),
            .I(N__16139));
    Glb2LocalMux I__2317 (
            .O(N__16204),
            .I(N__16139));
    Glb2LocalMux I__2316 (
            .O(N__16201),
            .I(N__16139));
    Glb2LocalMux I__2315 (
            .O(N__16198),
            .I(N__16139));
    Glb2LocalMux I__2314 (
            .O(N__16195),
            .I(N__16139));
    Glb2LocalMux I__2313 (
            .O(N__16192),
            .I(N__16139));
    GlobalMux I__2312 (
            .O(N__16139),
            .I(N__16136));
    gio2CtrlBuf I__2311 (
            .O(N__16136),
            .I(bram_enable_g));
    InMux I__2310 (
            .O(N__16133),
            .I(N__16130));
    LocalMux I__2309 (
            .O(N__16130),
            .I(N__16127));
    Odrv4 I__2308 (
            .O(N__16127),
            .I(\processor_zipi8.flags_i.m104Z0Z_2 ));
    InMux I__2307 (
            .O(N__16124),
            .I(N__16120));
    InMux I__2306 (
            .O(N__16123),
            .I(N__16117));
    LocalMux I__2305 (
            .O(N__16120),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6 ));
    LocalMux I__2304 (
            .O(N__16117),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6 ));
    InMux I__2303 (
            .O(N__16112),
            .I(N__16108));
    InMux I__2302 (
            .O(N__16111),
            .I(N__16105));
    LocalMux I__2301 (
            .O(N__16108),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6 ));
    LocalMux I__2300 (
            .O(N__16105),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6 ));
    CascadeMux I__2299 (
            .O(N__16100),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_6_cascade_ ));
    InMux I__2298 (
            .O(N__16097),
            .I(N__16094));
    LocalMux I__2297 (
            .O(N__16094),
            .I(N__16090));
    InMux I__2296 (
            .O(N__16093),
            .I(N__16087));
    Span4Mux_h I__2295 (
            .O(N__16090),
            .I(N__16082));
    LocalMux I__2294 (
            .O(N__16087),
            .I(N__16082));
    Odrv4 I__2293 (
            .O(N__16082),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_6 ));
    CascadeMux I__2292 (
            .O(N__16079),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI44F42_6_cascade_ ));
    CascadeMux I__2291 (
            .O(N__16076),
            .I(\processor_zipi8.decode4_strobes_enables_i.flag_enable_type_1_cascade_ ));
    InMux I__2290 (
            .O(N__16073),
            .I(N__16070));
    LocalMux I__2289 (
            .O(N__16070),
            .I(N__16067));
    Odrv12 I__2288 (
            .O(N__16067),
            .I(\processor_zipi8.shift_rotate_result_2 ));
    InMux I__2287 (
            .O(N__16064),
            .I(N__16061));
    LocalMux I__2286 (
            .O(N__16061),
            .I(N__16058));
    Span4Mux_v I__2285 (
            .O(N__16058),
            .I(N__16055));
    Odrv4 I__2284 (
            .O(N__16055),
            .I(\processor_zipi8.spm_data_2 ));
    CascadeMux I__2283 (
            .O(N__16052),
            .I(\processor_zipi8.register_bank_control_i.un31_regbank_type_3_cascade_ ));
    InMux I__2282 (
            .O(N__16049),
            .I(N__16046));
    LocalMux I__2281 (
            .O(N__16046),
            .I(N__16043));
    Odrv12 I__2280 (
            .O(N__16043),
            .I(\processor_zipi8.register_bank_control_i.un31_regbank_type ));
    InMux I__2279 (
            .O(N__16040),
            .I(N__16037));
    LocalMux I__2278 (
            .O(N__16037),
            .I(N__16034));
    Odrv12 I__2277 (
            .O(N__16034),
            .I(\processor_zipi8.shift_rotate_result_0 ));
    InMux I__2276 (
            .O(N__16031),
            .I(N__16028));
    LocalMux I__2275 (
            .O(N__16028),
            .I(N__16025));
    Span4Mux_v I__2274 (
            .O(N__16025),
            .I(N__16022));
    Span4Mux_v I__2273 (
            .O(N__16022),
            .I(N__16019));
    Odrv4 I__2272 (
            .O(N__16019),
            .I(\processor_zipi8.spm_data_0 ));
    CascadeMux I__2271 (
            .O(N__16016),
            .I(\processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_0_cascade_ ));
    InMux I__2270 (
            .O(N__16013),
            .I(N__16007));
    InMux I__2269 (
            .O(N__16012),
            .I(N__16007));
    LocalMux I__2268 (
            .O(N__16007),
            .I(N__16004));
    Span4Mux_v I__2267 (
            .O(N__16004),
            .I(N__16001));
    Odrv4 I__2266 (
            .O(N__16001),
            .I(\processor_zipi8.pc_mode_2_0_0 ));
    InMux I__2265 (
            .O(N__15998),
            .I(N__15995));
    LocalMux I__2264 (
            .O(N__15995),
            .I(N__15992));
    Odrv12 I__2263 (
            .O(N__15992),
            .I(\processor_zipi8.pc_vector_2 ));
    InMux I__2262 (
            .O(N__15989),
            .I(N__15986));
    LocalMux I__2261 (
            .O(N__15986),
            .I(N__15983));
    Odrv4 I__2260 (
            .O(N__15983),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_2 ));
    CascadeMux I__2259 (
            .O(N__15980),
            .I(N__15977));
    InMux I__2258 (
            .O(N__15977),
            .I(N__15971));
    InMux I__2257 (
            .O(N__15976),
            .I(N__15971));
    LocalMux I__2256 (
            .O(N__15971),
            .I(N__15967));
    InMux I__2255 (
            .O(N__15970),
            .I(N__15964));
    Odrv4 I__2254 (
            .O(N__15967),
            .I(\processor_zipi8.program_counter_i.half_pc_0_2 ));
    LocalMux I__2253 (
            .O(N__15964),
            .I(\processor_zipi8.program_counter_i.half_pc_0_2 ));
    InMux I__2252 (
            .O(N__15959),
            .I(N__15949));
    InMux I__2251 (
            .O(N__15958),
            .I(N__15949));
    InMux I__2250 (
            .O(N__15957),
            .I(N__15946));
    InMux I__2249 (
            .O(N__15956),
            .I(N__15941));
    InMux I__2248 (
            .O(N__15955),
            .I(N__15941));
    CascadeMux I__2247 (
            .O(N__15954),
            .I(N__15929));
    LocalMux I__2246 (
            .O(N__15949),
            .I(N__15921));
    LocalMux I__2245 (
            .O(N__15946),
            .I(N__15921));
    LocalMux I__2244 (
            .O(N__15941),
            .I(N__15918));
    InMux I__2243 (
            .O(N__15940),
            .I(N__15913));
    InMux I__2242 (
            .O(N__15939),
            .I(N__15913));
    InMux I__2241 (
            .O(N__15938),
            .I(N__15910));
    InMux I__2240 (
            .O(N__15937),
            .I(N__15903));
    InMux I__2239 (
            .O(N__15936),
            .I(N__15903));
    InMux I__2238 (
            .O(N__15935),
            .I(N__15903));
    InMux I__2237 (
            .O(N__15934),
            .I(N__15888));
    InMux I__2236 (
            .O(N__15933),
            .I(N__15888));
    InMux I__2235 (
            .O(N__15932),
            .I(N__15888));
    InMux I__2234 (
            .O(N__15929),
            .I(N__15888));
    InMux I__2233 (
            .O(N__15928),
            .I(N__15888));
    InMux I__2232 (
            .O(N__15927),
            .I(N__15888));
    InMux I__2231 (
            .O(N__15926),
            .I(N__15888));
    Span4Mux_v I__2230 (
            .O(N__15921),
            .I(N__15885));
    Span4Mux_h I__2229 (
            .O(N__15918),
            .I(N__15882));
    LocalMux I__2228 (
            .O(N__15913),
            .I(\processor_zipi8.program_counter_i.un3_half_pcZ0 ));
    LocalMux I__2227 (
            .O(N__15910),
            .I(\processor_zipi8.program_counter_i.un3_half_pcZ0 ));
    LocalMux I__2226 (
            .O(N__15903),
            .I(\processor_zipi8.program_counter_i.un3_half_pcZ0 ));
    LocalMux I__2225 (
            .O(N__15888),
            .I(\processor_zipi8.program_counter_i.un3_half_pcZ0 ));
    Odrv4 I__2224 (
            .O(N__15885),
            .I(\processor_zipi8.program_counter_i.un3_half_pcZ0 ));
    Odrv4 I__2223 (
            .O(N__15882),
            .I(\processor_zipi8.program_counter_i.un3_half_pcZ0 ));
    InMux I__2222 (
            .O(N__15869),
            .I(N__15866));
    LocalMux I__2221 (
            .O(N__15866),
            .I(N__15862));
    InMux I__2220 (
            .O(N__15865),
            .I(N__15859));
    Odrv4 I__2219 (
            .O(N__15862),
            .I(\processor_zipi8.program_counter_i.half_pc_0_3 ));
    LocalMux I__2218 (
            .O(N__15859),
            .I(\processor_zipi8.program_counter_i.half_pc_0_3 ));
    CascadeMux I__2217 (
            .O(N__15854),
            .I(\processor_zipi8.un16_alu_mux_sel_value_cascade_ ));
    InMux I__2216 (
            .O(N__15851),
            .I(N__15848));
    LocalMux I__2215 (
            .O(N__15848),
            .I(\processor_zipi8.decode4_strobes_enables_i.un23_flag_enable_type ));
    CascadeMux I__2214 (
            .O(N__15845),
            .I(\processor_zipi8.pc_vector_0_cascade_ ));
    InMux I__2213 (
            .O(N__15842),
            .I(N__15836));
    InMux I__2212 (
            .O(N__15841),
            .I(N__15836));
    LocalMux I__2211 (
            .O(N__15836),
            .I(N__15833));
    Span4Mux_h I__2210 (
            .O(N__15833),
            .I(N__15830));
    Odrv4 I__2209 (
            .O(N__15830),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_0 ));
    InMux I__2208 (
            .O(N__15827),
            .I(N__15823));
    CascadeMux I__2207 (
            .O(N__15826),
            .I(N__15820));
    LocalMux I__2206 (
            .O(N__15823),
            .I(N__15817));
    InMux I__2205 (
            .O(N__15820),
            .I(N__15814));
    Span4Mux_s3_h I__2204 (
            .O(N__15817),
            .I(N__15811));
    LocalMux I__2203 (
            .O(N__15814),
            .I(N__15808));
    Odrv4 I__2202 (
            .O(N__15811),
            .I(\processor_zipi8.flags_i.i14_mux ));
    Odrv12 I__2201 (
            .O(N__15808),
            .I(\processor_zipi8.flags_i.i14_mux ));
    InMux I__2200 (
            .O(N__15803),
            .I(N__15799));
    InMux I__2199 (
            .O(N__15802),
            .I(N__15796));
    LocalMux I__2198 (
            .O(N__15799),
            .I(N__15793));
    LocalMux I__2197 (
            .O(N__15796),
            .I(N__15790));
    Span4Mux_v I__2196 (
            .O(N__15793),
            .I(N__15787));
    Span4Mux_h I__2195 (
            .O(N__15790),
            .I(N__15784));
    Odrv4 I__2194 (
            .O(N__15787),
            .I(\processor_zipi8.flags_i.i14_mux_0 ));
    Odrv4 I__2193 (
            .O(N__15784),
            .I(\processor_zipi8.flags_i.i14_mux_0 ));
    CascadeMux I__2192 (
            .O(N__15779),
            .I(N__15776));
    InMux I__2191 (
            .O(N__15776),
            .I(N__15773));
    LocalMux I__2190 (
            .O(N__15773),
            .I(N__15770));
    Odrv4 I__2189 (
            .O(N__15770),
            .I(\processor_zipi8.zero_flag_RNIC4FP9 ));
    CEMux I__2188 (
            .O(N__15767),
            .I(N__15764));
    LocalMux I__2187 (
            .O(N__15764),
            .I(N__15759));
    CEMux I__2186 (
            .O(N__15763),
            .I(N__15755));
    CEMux I__2185 (
            .O(N__15762),
            .I(N__15752));
    Span4Mux_v I__2184 (
            .O(N__15759),
            .I(N__15749));
    CEMux I__2183 (
            .O(N__15758),
            .I(N__15746));
    LocalMux I__2182 (
            .O(N__15755),
            .I(N__15743));
    LocalMux I__2181 (
            .O(N__15752),
            .I(N__15740));
    Span4Mux_s1_h I__2180 (
            .O(N__15749),
            .I(N__15737));
    LocalMux I__2179 (
            .O(N__15746),
            .I(N__15734));
    Span4Mux_s2_h I__2178 (
            .O(N__15743),
            .I(N__15729));
    Span4Mux_s2_h I__2177 (
            .O(N__15740),
            .I(N__15729));
    Odrv4 I__2176 (
            .O(N__15737),
            .I(\processor_zipi8.program_counter_i.t_state_0_1 ));
    Odrv4 I__2175 (
            .O(N__15734),
            .I(\processor_zipi8.program_counter_i.t_state_0_1 ));
    Odrv4 I__2174 (
            .O(N__15729),
            .I(\processor_zipi8.program_counter_i.t_state_0_1 ));
    CascadeMux I__2173 (
            .O(N__15722),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_1_cascade_ ));
    CascadeMux I__2172 (
            .O(N__15719),
            .I(\processor_zipi8.program_counter_i.half_pc_0_1_cascade_ ));
    CascadeMux I__2171 (
            .O(N__15716),
            .I(N__15712));
    CascadeMux I__2170 (
            .O(N__15715),
            .I(N__15709));
    CascadeBuf I__2169 (
            .O(N__15712),
            .I(N__15706));
    CascadeBuf I__2168 (
            .O(N__15709),
            .I(N__15703));
    CascadeMux I__2167 (
            .O(N__15706),
            .I(N__15700));
    CascadeMux I__2166 (
            .O(N__15703),
            .I(N__15697));
    CascadeBuf I__2165 (
            .O(N__15700),
            .I(N__15694));
    CascadeBuf I__2164 (
            .O(N__15697),
            .I(N__15691));
    CascadeMux I__2163 (
            .O(N__15694),
            .I(N__15688));
    CascadeMux I__2162 (
            .O(N__15691),
            .I(N__15685));
    CascadeBuf I__2161 (
            .O(N__15688),
            .I(N__15682));
    CascadeBuf I__2160 (
            .O(N__15685),
            .I(N__15679));
    CascadeMux I__2159 (
            .O(N__15682),
            .I(N__15676));
    CascadeMux I__2158 (
            .O(N__15679),
            .I(N__15673));
    CascadeBuf I__2157 (
            .O(N__15676),
            .I(N__15670));
    CascadeBuf I__2156 (
            .O(N__15673),
            .I(N__15667));
    CascadeMux I__2155 (
            .O(N__15670),
            .I(N__15664));
    CascadeMux I__2154 (
            .O(N__15667),
            .I(N__15661));
    CascadeBuf I__2153 (
            .O(N__15664),
            .I(N__15658));
    CascadeBuf I__2152 (
            .O(N__15661),
            .I(N__15655));
    CascadeMux I__2151 (
            .O(N__15658),
            .I(N__15652));
    CascadeMux I__2150 (
            .O(N__15655),
            .I(N__15649));
    CascadeBuf I__2149 (
            .O(N__15652),
            .I(N__15646));
    CascadeBuf I__2148 (
            .O(N__15649),
            .I(N__15643));
    CascadeMux I__2147 (
            .O(N__15646),
            .I(N__15640));
    CascadeMux I__2146 (
            .O(N__15643),
            .I(N__15637));
    CascadeBuf I__2145 (
            .O(N__15640),
            .I(N__15634));
    CascadeBuf I__2144 (
            .O(N__15637),
            .I(N__15631));
    CascadeMux I__2143 (
            .O(N__15634),
            .I(N__15627));
    CascadeMux I__2142 (
            .O(N__15631),
            .I(N__15624));
    InMux I__2141 (
            .O(N__15630),
            .I(N__15621));
    InMux I__2140 (
            .O(N__15627),
            .I(N__15618));
    InMux I__2139 (
            .O(N__15624),
            .I(N__15615));
    LocalMux I__2138 (
            .O(N__15621),
            .I(N__15612));
    LocalMux I__2137 (
            .O(N__15618),
            .I(N__15606));
    LocalMux I__2136 (
            .O(N__15615),
            .I(N__15603));
    Span4Mux_v I__2135 (
            .O(N__15612),
            .I(N__15599));
    CascadeMux I__2134 (
            .O(N__15611),
            .I(N__15596));
    CascadeMux I__2133 (
            .O(N__15610),
            .I(N__15593));
    CascadeMux I__2132 (
            .O(N__15609),
            .I(N__15590));
    Span4Mux_v I__2131 (
            .O(N__15606),
            .I(N__15587));
    Span4Mux_s3_h I__2130 (
            .O(N__15603),
            .I(N__15584));
    InMux I__2129 (
            .O(N__15602),
            .I(N__15581));
    Sp12to4 I__2128 (
            .O(N__15599),
            .I(N__15578));
    InMux I__2127 (
            .O(N__15596),
            .I(N__15575));
    InMux I__2126 (
            .O(N__15593),
            .I(N__15572));
    InMux I__2125 (
            .O(N__15590),
            .I(N__15569));
    Span4Mux_h I__2124 (
            .O(N__15587),
            .I(N__15566));
    Span4Mux_h I__2123 (
            .O(N__15584),
            .I(N__15563));
    LocalMux I__2122 (
            .O(N__15581),
            .I(address_1));
    Odrv12 I__2121 (
            .O(N__15578),
            .I(address_1));
    LocalMux I__2120 (
            .O(N__15575),
            .I(address_1));
    LocalMux I__2119 (
            .O(N__15572),
            .I(address_1));
    LocalMux I__2118 (
            .O(N__15569),
            .I(address_1));
    Odrv4 I__2117 (
            .O(N__15566),
            .I(address_1));
    Odrv4 I__2116 (
            .O(N__15563),
            .I(address_1));
    InMux I__2115 (
            .O(N__15548),
            .I(N__15545));
    LocalMux I__2114 (
            .O(N__15545),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0 ));
    CascadeMux I__2113 (
            .O(N__15542),
            .I(N__15538));
    CascadeMux I__2112 (
            .O(N__15541),
            .I(N__15535));
    CascadeBuf I__2111 (
            .O(N__15538),
            .I(N__15532));
    CascadeBuf I__2110 (
            .O(N__15535),
            .I(N__15529));
    CascadeMux I__2109 (
            .O(N__15532),
            .I(N__15526));
    CascadeMux I__2108 (
            .O(N__15529),
            .I(N__15523));
    CascadeBuf I__2107 (
            .O(N__15526),
            .I(N__15520));
    CascadeBuf I__2106 (
            .O(N__15523),
            .I(N__15517));
    CascadeMux I__2105 (
            .O(N__15520),
            .I(N__15514));
    CascadeMux I__2104 (
            .O(N__15517),
            .I(N__15511));
    CascadeBuf I__2103 (
            .O(N__15514),
            .I(N__15508));
    CascadeBuf I__2102 (
            .O(N__15511),
            .I(N__15505));
    CascadeMux I__2101 (
            .O(N__15508),
            .I(N__15502));
    CascadeMux I__2100 (
            .O(N__15505),
            .I(N__15499));
    CascadeBuf I__2099 (
            .O(N__15502),
            .I(N__15496));
    CascadeBuf I__2098 (
            .O(N__15499),
            .I(N__15493));
    CascadeMux I__2097 (
            .O(N__15496),
            .I(N__15490));
    CascadeMux I__2096 (
            .O(N__15493),
            .I(N__15487));
    CascadeBuf I__2095 (
            .O(N__15490),
            .I(N__15484));
    CascadeBuf I__2094 (
            .O(N__15487),
            .I(N__15481));
    CascadeMux I__2093 (
            .O(N__15484),
            .I(N__15478));
    CascadeMux I__2092 (
            .O(N__15481),
            .I(N__15475));
    CascadeBuf I__2091 (
            .O(N__15478),
            .I(N__15472));
    CascadeBuf I__2090 (
            .O(N__15475),
            .I(N__15469));
    CascadeMux I__2089 (
            .O(N__15472),
            .I(N__15466));
    CascadeMux I__2088 (
            .O(N__15469),
            .I(N__15463));
    CascadeBuf I__2087 (
            .O(N__15466),
            .I(N__15460));
    CascadeBuf I__2086 (
            .O(N__15463),
            .I(N__15457));
    CascadeMux I__2085 (
            .O(N__15460),
            .I(N__15454));
    CascadeMux I__2084 (
            .O(N__15457),
            .I(N__15451));
    InMux I__2083 (
            .O(N__15454),
            .I(N__15445));
    InMux I__2082 (
            .O(N__15451),
            .I(N__15442));
    InMux I__2081 (
            .O(N__15450),
            .I(N__15438));
    InMux I__2080 (
            .O(N__15449),
            .I(N__15434));
    CascadeMux I__2079 (
            .O(N__15448),
            .I(N__15431));
    LocalMux I__2078 (
            .O(N__15445),
            .I(N__15426));
    LocalMux I__2077 (
            .O(N__15442),
            .I(N__15426));
    InMux I__2076 (
            .O(N__15441),
            .I(N__15423));
    LocalMux I__2075 (
            .O(N__15438),
            .I(N__15420));
    CascadeMux I__2074 (
            .O(N__15437),
            .I(N__15417));
    LocalMux I__2073 (
            .O(N__15434),
            .I(N__15414));
    InMux I__2072 (
            .O(N__15431),
            .I(N__15411));
    Span4Mux_v I__2071 (
            .O(N__15426),
            .I(N__15408));
    LocalMux I__2070 (
            .O(N__15423),
            .I(N__15403));
    Span4Mux_v I__2069 (
            .O(N__15420),
            .I(N__15403));
    InMux I__2068 (
            .O(N__15417),
            .I(N__15400));
    Span4Mux_v I__2067 (
            .O(N__15414),
            .I(N__15393));
    LocalMux I__2066 (
            .O(N__15411),
            .I(N__15393));
    Span4Mux_h I__2065 (
            .O(N__15408),
            .I(N__15393));
    Odrv4 I__2064 (
            .O(N__15403),
            .I(address_0));
    LocalMux I__2063 (
            .O(N__15400),
            .I(address_0));
    Odrv4 I__2062 (
            .O(N__15393),
            .I(address_0));
    CascadeMux I__2061 (
            .O(N__15386),
            .I(N__15383));
    InMux I__2060 (
            .O(N__15383),
            .I(N__15380));
    LocalMux I__2059 (
            .O(N__15380),
            .I(N__15377));
    Span4Mux_s3_h I__2058 (
            .O(N__15377),
            .I(N__15374));
    Odrv4 I__2057 (
            .O(N__15374),
            .I(\processor_zipi8.zero_flag_RNIL8RB5 ));
    InMux I__2056 (
            .O(N__15371),
            .I(N__15364));
    InMux I__2055 (
            .O(N__15370),
            .I(N__15364));
    CascadeMux I__2054 (
            .O(N__15369),
            .I(N__15361));
    LocalMux I__2053 (
            .O(N__15364),
            .I(N__15358));
    InMux I__2052 (
            .O(N__15361),
            .I(N__15355));
    Odrv4 I__2051 (
            .O(N__15358),
            .I(\processor_zipi8.program_counter_i.half_pc_0_1 ));
    LocalMux I__2050 (
            .O(N__15355),
            .I(\processor_zipi8.program_counter_i.half_pc_0_1 ));
    InMux I__2049 (
            .O(N__15350),
            .I(N__15342));
    InMux I__2048 (
            .O(N__15349),
            .I(N__15342));
    InMux I__2047 (
            .O(N__15348),
            .I(N__15337));
    InMux I__2046 (
            .O(N__15347),
            .I(N__15337));
    LocalMux I__2045 (
            .O(N__15342),
            .I(\processor_zipi8.program_counter_i.carry_pc_4_0 ));
    LocalMux I__2044 (
            .O(N__15337),
            .I(\processor_zipi8.program_counter_i.carry_pc_4_0 ));
    InMux I__2043 (
            .O(N__15332),
            .I(N__15326));
    InMux I__2042 (
            .O(N__15331),
            .I(N__15326));
    LocalMux I__2041 (
            .O(N__15326),
            .I(N__15323));
    Odrv4 I__2040 (
            .O(N__15323),
            .I(\processor_zipi8.program_counter_i.carry_pc_22_3 ));
    CascadeMux I__2039 (
            .O(N__15320),
            .I(N__15317));
    CascadeBuf I__2038 (
            .O(N__15317),
            .I(N__15314));
    CascadeMux I__2037 (
            .O(N__15314),
            .I(N__15310));
    CascadeMux I__2036 (
            .O(N__15313),
            .I(N__15307));
    CascadeBuf I__2035 (
            .O(N__15310),
            .I(N__15304));
    CascadeBuf I__2034 (
            .O(N__15307),
            .I(N__15301));
    CascadeMux I__2033 (
            .O(N__15304),
            .I(N__15298));
    CascadeMux I__2032 (
            .O(N__15301),
            .I(N__15295));
    CascadeBuf I__2031 (
            .O(N__15298),
            .I(N__15292));
    CascadeBuf I__2030 (
            .O(N__15295),
            .I(N__15289));
    CascadeMux I__2029 (
            .O(N__15292),
            .I(N__15286));
    CascadeMux I__2028 (
            .O(N__15289),
            .I(N__15283));
    CascadeBuf I__2027 (
            .O(N__15286),
            .I(N__15280));
    CascadeBuf I__2026 (
            .O(N__15283),
            .I(N__15277));
    CascadeMux I__2025 (
            .O(N__15280),
            .I(N__15274));
    CascadeMux I__2024 (
            .O(N__15277),
            .I(N__15271));
    CascadeBuf I__2023 (
            .O(N__15274),
            .I(N__15268));
    CascadeBuf I__2022 (
            .O(N__15271),
            .I(N__15265));
    CascadeMux I__2021 (
            .O(N__15268),
            .I(N__15262));
    CascadeMux I__2020 (
            .O(N__15265),
            .I(N__15259));
    CascadeBuf I__2019 (
            .O(N__15262),
            .I(N__15256));
    CascadeBuf I__2018 (
            .O(N__15259),
            .I(N__15253));
    CascadeMux I__2017 (
            .O(N__15256),
            .I(N__15250));
    CascadeMux I__2016 (
            .O(N__15253),
            .I(N__15247));
    CascadeBuf I__2015 (
            .O(N__15250),
            .I(N__15244));
    CascadeBuf I__2014 (
            .O(N__15247),
            .I(N__15241));
    CascadeMux I__2013 (
            .O(N__15244),
            .I(N__15238));
    CascadeMux I__2012 (
            .O(N__15241),
            .I(N__15235));
    InMux I__2011 (
            .O(N__15238),
            .I(N__15231));
    CascadeBuf I__2010 (
            .O(N__15235),
            .I(N__15228));
    CascadeMux I__2009 (
            .O(N__15234),
            .I(N__15224));
    LocalMux I__2008 (
            .O(N__15231),
            .I(N__15221));
    CascadeMux I__2007 (
            .O(N__15228),
            .I(N__15218));
    InMux I__2006 (
            .O(N__15227),
            .I(N__15215));
    InMux I__2005 (
            .O(N__15224),
            .I(N__15211));
    Span4Mux_s1_v I__2004 (
            .O(N__15221),
            .I(N__15208));
    InMux I__2003 (
            .O(N__15218),
            .I(N__15205));
    LocalMux I__2002 (
            .O(N__15215),
            .I(N__15201));
    CascadeMux I__2001 (
            .O(N__15214),
            .I(N__15198));
    LocalMux I__2000 (
            .O(N__15211),
            .I(N__15195));
    Sp12to4 I__1999 (
            .O(N__15208),
            .I(N__15190));
    LocalMux I__1998 (
            .O(N__15205),
            .I(N__15190));
    InMux I__1997 (
            .O(N__15204),
            .I(N__15187));
    Span4Mux_s3_h I__1996 (
            .O(N__15201),
            .I(N__15184));
    InMux I__1995 (
            .O(N__15198),
            .I(N__15181));
    Sp12to4 I__1994 (
            .O(N__15195),
            .I(N__15176));
    Span12Mux_s8_h I__1993 (
            .O(N__15190),
            .I(N__15176));
    LocalMux I__1992 (
            .O(N__15187),
            .I(address_2));
    Odrv4 I__1991 (
            .O(N__15184),
            .I(address_2));
    LocalMux I__1990 (
            .O(N__15181),
            .I(address_2));
    Odrv12 I__1989 (
            .O(N__15176),
            .I(address_2));
    CascadeMux I__1988 (
            .O(N__15167),
            .I(N__15162));
    CascadeMux I__1987 (
            .O(N__15166),
            .I(N__15159));
    InMux I__1986 (
            .O(N__15165),
            .I(N__15154));
    InMux I__1985 (
            .O(N__15162),
            .I(N__15151));
    InMux I__1984 (
            .O(N__15159),
            .I(N__15148));
    CascadeMux I__1983 (
            .O(N__15158),
            .I(N__15145));
    InMux I__1982 (
            .O(N__15157),
            .I(N__15141));
    LocalMux I__1981 (
            .O(N__15154),
            .I(N__15136));
    LocalMux I__1980 (
            .O(N__15151),
            .I(N__15136));
    LocalMux I__1979 (
            .O(N__15148),
            .I(N__15133));
    InMux I__1978 (
            .O(N__15145),
            .I(N__15128));
    InMux I__1977 (
            .O(N__15144),
            .I(N__15128));
    LocalMux I__1976 (
            .O(N__15141),
            .I(N__15125));
    Span4Mux_s2_v I__1975 (
            .O(N__15136),
            .I(N__15122));
    Odrv4 I__1974 (
            .O(N__15133),
            .I(\processor_zipi8.stack_pointer_4 ));
    LocalMux I__1973 (
            .O(N__15128),
            .I(\processor_zipi8.stack_pointer_4 ));
    Odrv4 I__1972 (
            .O(N__15125),
            .I(\processor_zipi8.stack_pointer_4 ));
    Odrv4 I__1971 (
            .O(N__15122),
            .I(\processor_zipi8.stack_pointer_4 ));
    CascadeMux I__1970 (
            .O(N__15113),
            .I(N__15110));
    InMux I__1969 (
            .O(N__15110),
            .I(N__15106));
    InMux I__1968 (
            .O(N__15109),
            .I(N__15103));
    LocalMux I__1967 (
            .O(N__15106),
            .I(N__15097));
    LocalMux I__1966 (
            .O(N__15103),
            .I(N__15097));
    InMux I__1965 (
            .O(N__15102),
            .I(N__15094));
    Span4Mux_h I__1964 (
            .O(N__15097),
            .I(N__15091));
    LocalMux I__1963 (
            .O(N__15094),
            .I(N__15088));
    Odrv4 I__1962 (
            .O(N__15091),
            .I(\processor_zipi8.flags_i.N_34 ));
    Odrv4 I__1961 (
            .O(N__15088),
            .I(\processor_zipi8.flags_i.N_34 ));
    CascadeMux I__1960 (
            .O(N__15083),
            .I(\processor_zipi8.port_id_0_cascade_ ));
    InMux I__1959 (
            .O(N__15080),
            .I(N__15077));
    LocalMux I__1958 (
            .O(N__15077),
            .I(N__15074));
    Span4Mux_v I__1957 (
            .O(N__15074),
            .I(N__15071));
    Odrv4 I__1956 (
            .O(N__15071),
            .I(\processor_zipi8.stack_memory_0 ));
    InMux I__1955 (
            .O(N__15068),
            .I(N__15065));
    LocalMux I__1954 (
            .O(N__15065),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_0 ));
    CascadeMux I__1953 (
            .O(N__15062),
            .I(N__15059));
    InMux I__1952 (
            .O(N__15059),
            .I(N__15056));
    LocalMux I__1951 (
            .O(N__15056),
            .I(N__15053));
    Odrv4 I__1950 (
            .O(N__15053),
            .I(\processor_zipi8.pc_vector_0 ));
    CascadeMux I__1949 (
            .O(N__15050),
            .I(N__15046));
    CascadeMux I__1948 (
            .O(N__15049),
            .I(N__15042));
    InMux I__1947 (
            .O(N__15046),
            .I(N__15039));
    CascadeMux I__1946 (
            .O(N__15045),
            .I(N__15036));
    InMux I__1945 (
            .O(N__15042),
            .I(N__15031));
    LocalMux I__1944 (
            .O(N__15039),
            .I(N__15028));
    InMux I__1943 (
            .O(N__15036),
            .I(N__15025));
    InMux I__1942 (
            .O(N__15035),
            .I(N__15020));
    InMux I__1941 (
            .O(N__15034),
            .I(N__15020));
    LocalMux I__1940 (
            .O(N__15031),
            .I(\processor_zipi8.port_id_2 ));
    Odrv4 I__1939 (
            .O(N__15028),
            .I(\processor_zipi8.port_id_2 ));
    LocalMux I__1938 (
            .O(N__15025),
            .I(\processor_zipi8.port_id_2 ));
    LocalMux I__1937 (
            .O(N__15020),
            .I(\processor_zipi8.port_id_2 ));
    InMux I__1936 (
            .O(N__15011),
            .I(N__15008));
    LocalMux I__1935 (
            .O(N__15008),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_2 ));
    InMux I__1934 (
            .O(N__15005),
            .I(N__15002));
    LocalMux I__1933 (
            .O(N__15002),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_2 ));
    CascadeMux I__1932 (
            .O(N__14999),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_2_cascade_ ));
    InMux I__1931 (
            .O(N__14996),
            .I(N__14993));
    LocalMux I__1930 (
            .O(N__14993),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_2 ));
    InMux I__1929 (
            .O(N__14990),
            .I(N__14987));
    LocalMux I__1928 (
            .O(N__14987),
            .I(N__14984));
    Span4Mux_h I__1927 (
            .O(N__14984),
            .I(N__14981));
    Odrv4 I__1926 (
            .O(N__14981),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_2 ));
    CascadeMux I__1925 (
            .O(N__14978),
            .I(\processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_0_cascade_ ));
    CascadeMux I__1924 (
            .O(N__14975),
            .I(N__14970));
    InMux I__1923 (
            .O(N__14974),
            .I(N__14961));
    InMux I__1922 (
            .O(N__14973),
            .I(N__14961));
    InMux I__1921 (
            .O(N__14970),
            .I(N__14961));
    InMux I__1920 (
            .O(N__14969),
            .I(N__14958));
    InMux I__1919 (
            .O(N__14968),
            .I(N__14955));
    LocalMux I__1918 (
            .O(N__14961),
            .I(N__14948));
    LocalMux I__1917 (
            .O(N__14958),
            .I(N__14948));
    LocalMux I__1916 (
            .O(N__14955),
            .I(N__14948));
    Span4Mux_v I__1915 (
            .O(N__14948),
            .I(N__14945));
    Span4Mux_v I__1914 (
            .O(N__14945),
            .I(N__14942));
    Span4Mux_h I__1913 (
            .O(N__14942),
            .I(N__14939));
    Odrv4 I__1912 (
            .O(N__14939),
            .I(instruction_2));
    CascadeMux I__1911 (
            .O(N__14936),
            .I(\processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_1_cascade_ ));
    InMux I__1910 (
            .O(N__14933),
            .I(N__14927));
    InMux I__1909 (
            .O(N__14932),
            .I(N__14927));
    LocalMux I__1908 (
            .O(N__14927),
            .I(N__14924));
    Odrv4 I__1907 (
            .O(N__14924),
            .I(\processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_0 ));
    InMux I__1906 (
            .O(N__14921),
            .I(N__14918));
    LocalMux I__1905 (
            .O(N__14918),
            .I(N__14915));
    Odrv12 I__1904 (
            .O(N__14915),
            .I(\processor_zipi8.shift_rotate_result_6 ));
    InMux I__1903 (
            .O(N__14912),
            .I(N__14909));
    LocalMux I__1902 (
            .O(N__14909),
            .I(N__14906));
    Span4Mux_s3_h I__1901 (
            .O(N__14906),
            .I(N__14903));
    Odrv4 I__1900 (
            .O(N__14903),
            .I(\processor_zipi8.shift_rotate_result_5 ));
    CascadeMux I__1899 (
            .O(N__14900),
            .I(\processor_zipi8.port_id_2_cascade_ ));
    CEMux I__1898 (
            .O(N__14897),
            .I(N__14894));
    LocalMux I__1897 (
            .O(N__14894),
            .I(N__14891));
    Span4Mux_s3_h I__1896 (
            .O(N__14891),
            .I(N__14888));
    Odrv4 I__1895 (
            .O(N__14888),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe11 ));
    CascadeMux I__1894 (
            .O(N__14885),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212_cascade_ ));
    InMux I__1893 (
            .O(N__14882),
            .I(N__14879));
    LocalMux I__1892 (
            .O(N__14879),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_0 ));
    CEMux I__1891 (
            .O(N__14876),
            .I(N__14873));
    LocalMux I__1890 (
            .O(N__14873),
            .I(N__14870));
    Span4Mux_s3_h I__1889 (
            .O(N__14870),
            .I(N__14867));
    Odrv4 I__1888 (
            .O(N__14867),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe8 ));
    CEMux I__1887 (
            .O(N__14864),
            .I(N__14860));
    CEMux I__1886 (
            .O(N__14863),
            .I(N__14857));
    LocalMux I__1885 (
            .O(N__14860),
            .I(N__14854));
    LocalMux I__1884 (
            .O(N__14857),
            .I(N__14851));
    Span4Mux_s1_v I__1883 (
            .O(N__14854),
            .I(N__14848));
    Span4Mux_s3_h I__1882 (
            .O(N__14851),
            .I(N__14845));
    Span4Mux_v I__1881 (
            .O(N__14848),
            .I(N__14842));
    Span4Mux_h I__1880 (
            .O(N__14845),
            .I(N__14839));
    Odrv4 I__1879 (
            .O(N__14842),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10 ));
    Odrv4 I__1878 (
            .O(N__14839),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10 ));
    CascadeMux I__1877 (
            .O(N__14834),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268_cascade_ ));
    InMux I__1876 (
            .O(N__14831),
            .I(N__14828));
    LocalMux I__1875 (
            .O(N__14828),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_6 ));
    InMux I__1874 (
            .O(N__14825),
            .I(N__14819));
    InMux I__1873 (
            .O(N__14824),
            .I(N__14819));
    LocalMux I__1872 (
            .O(N__14819),
            .I(N__14816));
    Span4Mux_h I__1871 (
            .O(N__14816),
            .I(N__14813));
    Odrv4 I__1870 (
            .O(N__14813),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_0 ));
    InMux I__1869 (
            .O(N__14810),
            .I(N__14804));
    InMux I__1868 (
            .O(N__14809),
            .I(N__14804));
    LocalMux I__1867 (
            .O(N__14804),
            .I(N__14801));
    Span4Mux_h I__1866 (
            .O(N__14801),
            .I(N__14798));
    Odrv4 I__1865 (
            .O(N__14798),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_0 ));
    CascadeMux I__1864 (
            .O(N__14795),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_0_cascade_ ));
    InMux I__1863 (
            .O(N__14792),
            .I(N__14786));
    InMux I__1862 (
            .O(N__14791),
            .I(N__14786));
    LocalMux I__1861 (
            .O(N__14786),
            .I(N__14783));
    Sp12to4 I__1860 (
            .O(N__14783),
            .I(N__14780));
    Odrv12 I__1859 (
            .O(N__14780),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_0 ));
    CascadeMux I__1858 (
            .O(N__14777),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_0_cascade_ ));
    InMux I__1857 (
            .O(N__14774),
            .I(N__14771));
    LocalMux I__1856 (
            .O(N__14771),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_0 ));
    CascadeMux I__1855 (
            .O(N__14768),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_0_cascade_ ));
    InMux I__1854 (
            .O(N__14765),
            .I(N__14762));
    LocalMux I__1853 (
            .O(N__14762),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_0 ));
    CascadeMux I__1852 (
            .O(N__14759),
            .I(\processor_zipi8.flags_i.m68_ns_1_cascade_ ));
    CascadeMux I__1851 (
            .O(N__14756),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_6_cascade_ ));
    InMux I__1850 (
            .O(N__14753),
            .I(N__14750));
    LocalMux I__1849 (
            .O(N__14750),
            .I(N__14747));
    Odrv4 I__1848 (
            .O(N__14747),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_6 ));
    InMux I__1847 (
            .O(N__14744),
            .I(N__14741));
    LocalMux I__1846 (
            .O(N__14741),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_6 ));
    CascadeMux I__1845 (
            .O(N__14738),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_6_cascade_ ));
    InMux I__1844 (
            .O(N__14735),
            .I(N__14732));
    LocalMux I__1843 (
            .O(N__14732),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_6 ));
    InMux I__1842 (
            .O(N__14729),
            .I(N__14726));
    LocalMux I__1841 (
            .O(N__14726),
            .I(N__14723));
    Span4Mux_h I__1840 (
            .O(N__14723),
            .I(N__14720));
    Odrv4 I__1839 (
            .O(N__14720),
            .I(\processor_zipi8.spm_data_6 ));
    CascadeMux I__1838 (
            .O(N__14717),
            .I(\processor_zipi8.flags_i.N_1235_cascade_ ));
    InMux I__1837 (
            .O(N__14714),
            .I(N__14711));
    LocalMux I__1836 (
            .O(N__14711),
            .I(\processor_zipi8.flags_i.zero_flag_RNI89VZ0Z91 ));
    CascadeMux I__1835 (
            .O(N__14708),
            .I(N__14705));
    InMux I__1834 (
            .O(N__14705),
            .I(N__14702));
    LocalMux I__1833 (
            .O(N__14702),
            .I(\processor_zipi8.flags_i.N_1239 ));
    InMux I__1832 (
            .O(N__14699),
            .I(N__14696));
    LocalMux I__1831 (
            .O(N__14696),
            .I(\processor_zipi8.flags_i.N_124_mux ));
    CascadeMux I__1830 (
            .O(N__14693),
            .I(\processor_zipi8.flags_i.N_1241_cascade_ ));
    CascadeMux I__1829 (
            .O(N__14690),
            .I(N__14687));
    InMux I__1828 (
            .O(N__14687),
            .I(N__14684));
    LocalMux I__1827 (
            .O(N__14684),
            .I(N__14681));
    Span4Mux_v I__1826 (
            .O(N__14681),
            .I(N__14678));
    Odrv4 I__1825 (
            .O(N__14678),
            .I(\processor_zipi8.zero_flag_RNIDS654 ));
    CascadeMux I__1824 (
            .O(N__14675),
            .I(N__14672));
    InMux I__1823 (
            .O(N__14672),
            .I(N__14669));
    LocalMux I__1822 (
            .O(N__14669),
            .I(N__14666));
    Span4Mux_h I__1821 (
            .O(N__14666),
            .I(N__14663));
    Span4Mux_v I__1820 (
            .O(N__14663),
            .I(N__14654));
    InMux I__1819 (
            .O(N__14662),
            .I(N__14651));
    InMux I__1818 (
            .O(N__14661),
            .I(N__14648));
    InMux I__1817 (
            .O(N__14660),
            .I(N__14643));
    InMux I__1816 (
            .O(N__14659),
            .I(N__14643));
    InMux I__1815 (
            .O(N__14658),
            .I(N__14640));
    InMux I__1814 (
            .O(N__14657),
            .I(N__14637));
    Odrv4 I__1813 (
            .O(N__14654),
            .I(\processor_zipi8.stack_pointer_1 ));
    LocalMux I__1812 (
            .O(N__14651),
            .I(\processor_zipi8.stack_pointer_1 ));
    LocalMux I__1811 (
            .O(N__14648),
            .I(\processor_zipi8.stack_pointer_1 ));
    LocalMux I__1810 (
            .O(N__14643),
            .I(\processor_zipi8.stack_pointer_1 ));
    LocalMux I__1809 (
            .O(N__14640),
            .I(\processor_zipi8.stack_pointer_1 ));
    LocalMux I__1808 (
            .O(N__14637),
            .I(\processor_zipi8.stack_pointer_1 ));
    CascadeMux I__1807 (
            .O(N__14624),
            .I(N__14621));
    InMux I__1806 (
            .O(N__14621),
            .I(N__14618));
    LocalMux I__1805 (
            .O(N__14618),
            .I(\processor_zipi8.flags_i.m75_amZ0 ));
    CascadeMux I__1804 (
            .O(N__14615),
            .I(\processor_zipi8.flags_i.m75_amZ0_cascade_ ));
    InMux I__1803 (
            .O(N__14612),
            .I(N__14606));
    InMux I__1802 (
            .O(N__14611),
            .I(N__14606));
    LocalMux I__1801 (
            .O(N__14606),
            .I(\processor_zipi8.flags_i.zero_flag_RNI3VCZ0Z94 ));
    CascadeMux I__1800 (
            .O(N__14603),
            .I(N__14600));
    InMux I__1799 (
            .O(N__14600),
            .I(N__14597));
    LocalMux I__1798 (
            .O(N__14597),
            .I(N__14594));
    Span4Mux_v I__1797 (
            .O(N__14594),
            .I(N__14591));
    Odrv4 I__1796 (
            .O(N__14591),
            .I(\processor_zipi8.zero_flag_RNI5GK75 ));
    InMux I__1795 (
            .O(N__14588),
            .I(N__14585));
    LocalMux I__1794 (
            .O(N__14585),
            .I(\processor_zipi8.flags_i.N_1241 ));
    CascadeMux I__1793 (
            .O(N__14582),
            .I(N__14579));
    InMux I__1792 (
            .O(N__14579),
            .I(N__14574));
    CascadeMux I__1791 (
            .O(N__14578),
            .I(N__14570));
    CascadeMux I__1790 (
            .O(N__14577),
            .I(N__14564));
    LocalMux I__1789 (
            .O(N__14574),
            .I(N__14561));
    CascadeMux I__1788 (
            .O(N__14573),
            .I(N__14556));
    InMux I__1787 (
            .O(N__14570),
            .I(N__14548));
    InMux I__1786 (
            .O(N__14569),
            .I(N__14548));
    InMux I__1785 (
            .O(N__14568),
            .I(N__14541));
    InMux I__1784 (
            .O(N__14567),
            .I(N__14541));
    InMux I__1783 (
            .O(N__14564),
            .I(N__14541));
    Span4Mux_v I__1782 (
            .O(N__14561),
            .I(N__14538));
    InMux I__1781 (
            .O(N__14560),
            .I(N__14533));
    InMux I__1780 (
            .O(N__14559),
            .I(N__14533));
    InMux I__1779 (
            .O(N__14556),
            .I(N__14530));
    InMux I__1778 (
            .O(N__14555),
            .I(N__14527));
    InMux I__1777 (
            .O(N__14554),
            .I(N__14524));
    InMux I__1776 (
            .O(N__14553),
            .I(N__14521));
    LocalMux I__1775 (
            .O(N__14548),
            .I(N__14516));
    LocalMux I__1774 (
            .O(N__14541),
            .I(N__14516));
    Odrv4 I__1773 (
            .O(N__14538),
            .I(\processor_zipi8.stack_pointer_0 ));
    LocalMux I__1772 (
            .O(N__14533),
            .I(\processor_zipi8.stack_pointer_0 ));
    LocalMux I__1771 (
            .O(N__14530),
            .I(\processor_zipi8.stack_pointer_0 ));
    LocalMux I__1770 (
            .O(N__14527),
            .I(\processor_zipi8.stack_pointer_0 ));
    LocalMux I__1769 (
            .O(N__14524),
            .I(\processor_zipi8.stack_pointer_0 ));
    LocalMux I__1768 (
            .O(N__14521),
            .I(\processor_zipi8.stack_pointer_0 ));
    Odrv4 I__1767 (
            .O(N__14516),
            .I(\processor_zipi8.stack_pointer_0 ));
    CascadeMux I__1766 (
            .O(N__14501),
            .I(N__14498));
    InMux I__1765 (
            .O(N__14498),
            .I(N__14495));
    LocalMux I__1764 (
            .O(N__14495),
            .I(N__14492));
    Span4Mux_v I__1763 (
            .O(N__14492),
            .I(N__14488));
    InMux I__1762 (
            .O(N__14491),
            .I(N__14481));
    Span4Mux_v I__1761 (
            .O(N__14488),
            .I(N__14478));
    InMux I__1760 (
            .O(N__14487),
            .I(N__14473));
    InMux I__1759 (
            .O(N__14486),
            .I(N__14473));
    InMux I__1758 (
            .O(N__14485),
            .I(N__14468));
    InMux I__1757 (
            .O(N__14484),
            .I(N__14468));
    LocalMux I__1756 (
            .O(N__14481),
            .I(N__14465));
    Odrv4 I__1755 (
            .O(N__14478),
            .I(\processor_zipi8.stack_pointer_2 ));
    LocalMux I__1754 (
            .O(N__14473),
            .I(\processor_zipi8.stack_pointer_2 ));
    LocalMux I__1753 (
            .O(N__14468),
            .I(\processor_zipi8.stack_pointer_2 ));
    Odrv4 I__1752 (
            .O(N__14465),
            .I(\processor_zipi8.stack_pointer_2 ));
    InMux I__1751 (
            .O(N__14456),
            .I(N__14449));
    InMux I__1750 (
            .O(N__14455),
            .I(N__14449));
    InMux I__1749 (
            .O(N__14454),
            .I(N__14446));
    LocalMux I__1748 (
            .O(N__14449),
            .I(\processor_zipi8.flags_i.N_54 ));
    LocalMux I__1747 (
            .O(N__14446),
            .I(\processor_zipi8.flags_i.N_54 ));
    CascadeMux I__1746 (
            .O(N__14441),
            .I(\processor_zipi8.flags_i.m91_amZ0_cascade_ ));
    CascadeMux I__1745 (
            .O(N__14438),
            .I(\processor_zipi8.flags_i.m25_ns_1_cascade_ ));
    CascadeMux I__1744 (
            .O(N__14435),
            .I(\processor_zipi8.flags_i.N_26_0_cascade_ ));
    InMux I__1743 (
            .O(N__14432),
            .I(N__14429));
    LocalMux I__1742 (
            .O(N__14429),
            .I(\processor_zipi8.flags_i.N_27_0 ));
    CascadeMux I__1741 (
            .O(N__14426),
            .I(\processor_zipi8.flags_i.m20_ns_1_cascade_ ));
    InMux I__1740 (
            .O(N__14423),
            .I(N__14420));
    LocalMux I__1739 (
            .O(N__14420),
            .I(\processor_zipi8.flags_i.N_21_0 ));
    InMux I__1738 (
            .O(N__14417),
            .I(N__14414));
    LocalMux I__1737 (
            .O(N__14414),
            .I(\processor_zipi8.program_counter_i.half_pc_0_10 ));
    InMux I__1736 (
            .O(N__14411),
            .I(N__14408));
    LocalMux I__1735 (
            .O(N__14408),
            .I(\processor_zipi8.program_counter_i.un431_half_pc ));
    CascadeMux I__1734 (
            .O(N__14405),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_11_cascade_ ));
    InMux I__1733 (
            .O(N__14402),
            .I(N__14399));
    LocalMux I__1732 (
            .O(N__14399),
            .I(N__14395));
    InMux I__1731 (
            .O(N__14398),
            .I(N__14392));
    Odrv4 I__1730 (
            .O(N__14395),
            .I(\processor_zipi8.address_11 ));
    LocalMux I__1729 (
            .O(N__14392),
            .I(\processor_zipi8.address_11 ));
    InMux I__1728 (
            .O(N__14387),
            .I(N__14384));
    LocalMux I__1727 (
            .O(N__14384),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_9 ));
    CascadeMux I__1726 (
            .O(N__14381),
            .I(N__14377));
    InMux I__1725 (
            .O(N__14380),
            .I(N__14374));
    InMux I__1724 (
            .O(N__14377),
            .I(N__14371));
    LocalMux I__1723 (
            .O(N__14374),
            .I(\processor_zipi8.pc_vector_9 ));
    LocalMux I__1722 (
            .O(N__14371),
            .I(\processor_zipi8.pc_vector_9 ));
    InMux I__1721 (
            .O(N__14366),
            .I(N__14362));
    InMux I__1720 (
            .O(N__14365),
            .I(N__14359));
    LocalMux I__1719 (
            .O(N__14362),
            .I(\processor_zipi8.program_counter_i.carry_pc_52_8 ));
    LocalMux I__1718 (
            .O(N__14359),
            .I(\processor_zipi8.program_counter_i.carry_pc_52_8 ));
    InMux I__1717 (
            .O(N__14354),
            .I(N__14350));
    InMux I__1716 (
            .O(N__14353),
            .I(N__14347));
    LocalMux I__1715 (
            .O(N__14350),
            .I(\processor_zipi8.program_counter_i.carry_pc_58_9 ));
    LocalMux I__1714 (
            .O(N__14347),
            .I(\processor_zipi8.program_counter_i.carry_pc_58_9 ));
    CascadeMux I__1713 (
            .O(N__14342),
            .I(N__14339));
    InMux I__1712 (
            .O(N__14339),
            .I(N__14336));
    LocalMux I__1711 (
            .O(N__14336),
            .I(\processor_zipi8.flags_i.m49_ns_1 ));
    CascadeMux I__1710 (
            .O(N__14333),
            .I(\processor_zipi8.flags_i.N_50_cascade_ ));
    CascadeMux I__1709 (
            .O(N__14330),
            .I(\processor_zipi8.flags_i.N_51_cascade_ ));
    InMux I__1708 (
            .O(N__14327),
            .I(N__14318));
    InMux I__1707 (
            .O(N__14326),
            .I(N__14318));
    InMux I__1706 (
            .O(N__14325),
            .I(N__14318));
    LocalMux I__1705 (
            .O(N__14318),
            .I(\processor_zipi8.flags_i.N_123_mux ));
    InMux I__1704 (
            .O(N__14315),
            .I(N__14312));
    LocalMux I__1703 (
            .O(N__14312),
            .I(\processor_zipi8.flags_i.N_45 ));
    CascadeMux I__1702 (
            .O(N__14309),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_4_cascade_ ));
    CascadeMux I__1701 (
            .O(N__14306),
            .I(\processor_zipi8.program_counter_i.carry_pc_28_4_cascade_ ));
    InMux I__1700 (
            .O(N__14303),
            .I(N__14300));
    LocalMux I__1699 (
            .O(N__14300),
            .I(\processor_zipi8.program_counter_i.carry_pc_34_5 ));
    CascadeMux I__1698 (
            .O(N__14297),
            .I(N__14294));
    InMux I__1697 (
            .O(N__14294),
            .I(N__14288));
    InMux I__1696 (
            .O(N__14293),
            .I(N__14288));
    LocalMux I__1695 (
            .O(N__14288),
            .I(N__14285));
    Span4Mux_s2_h I__1694 (
            .O(N__14285),
            .I(N__14282));
    Odrv4 I__1693 (
            .O(N__14282),
            .I(\processor_zipi8.pc_vector_6 ));
    CascadeMux I__1692 (
            .O(N__14279),
            .I(\processor_zipi8.program_counter_i.carry_pc_34_5_cascade_ ));
    InMux I__1691 (
            .O(N__14276),
            .I(N__14270));
    InMux I__1690 (
            .O(N__14275),
            .I(N__14270));
    LocalMux I__1689 (
            .O(N__14270),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_6 ));
    InMux I__1688 (
            .O(N__14267),
            .I(N__14264));
    LocalMux I__1687 (
            .O(N__14264),
            .I(\processor_zipi8.program_counter_i.carry_pc_40_6 ));
    CascadeMux I__1686 (
            .O(N__14261),
            .I(N__14257));
    InMux I__1685 (
            .O(N__14260),
            .I(N__14254));
    InMux I__1684 (
            .O(N__14257),
            .I(N__14251));
    LocalMux I__1683 (
            .O(N__14254),
            .I(N__14248));
    LocalMux I__1682 (
            .O(N__14251),
            .I(N__14245));
    Odrv4 I__1681 (
            .O(N__14248),
            .I(\processor_zipi8.pc_vector_7 ));
    Odrv12 I__1680 (
            .O(N__14245),
            .I(\processor_zipi8.pc_vector_7 ));
    CascadeMux I__1679 (
            .O(N__14240),
            .I(\processor_zipi8.program_counter_i.carry_pc_40_6_cascade_ ));
    InMux I__1678 (
            .O(N__14237),
            .I(N__14233));
    InMux I__1677 (
            .O(N__14236),
            .I(N__14230));
    LocalMux I__1676 (
            .O(N__14233),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_7 ));
    LocalMux I__1675 (
            .O(N__14230),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_7 ));
    CascadeMux I__1674 (
            .O(N__14225),
            .I(N__14222));
    CascadeBuf I__1673 (
            .O(N__14222),
            .I(N__14218));
    CascadeMux I__1672 (
            .O(N__14221),
            .I(N__14215));
    CascadeMux I__1671 (
            .O(N__14218),
            .I(N__14212));
    CascadeBuf I__1670 (
            .O(N__14215),
            .I(N__14209));
    CascadeBuf I__1669 (
            .O(N__14212),
            .I(N__14206));
    CascadeMux I__1668 (
            .O(N__14209),
            .I(N__14203));
    CascadeMux I__1667 (
            .O(N__14206),
            .I(N__14200));
    CascadeBuf I__1666 (
            .O(N__14203),
            .I(N__14197));
    CascadeBuf I__1665 (
            .O(N__14200),
            .I(N__14194));
    CascadeMux I__1664 (
            .O(N__14197),
            .I(N__14191));
    CascadeMux I__1663 (
            .O(N__14194),
            .I(N__14188));
    CascadeBuf I__1662 (
            .O(N__14191),
            .I(N__14185));
    CascadeBuf I__1661 (
            .O(N__14188),
            .I(N__14182));
    CascadeMux I__1660 (
            .O(N__14185),
            .I(N__14179));
    CascadeMux I__1659 (
            .O(N__14182),
            .I(N__14176));
    CascadeBuf I__1658 (
            .O(N__14179),
            .I(N__14173));
    CascadeBuf I__1657 (
            .O(N__14176),
            .I(N__14170));
    CascadeMux I__1656 (
            .O(N__14173),
            .I(N__14167));
    CascadeMux I__1655 (
            .O(N__14170),
            .I(N__14164));
    CascadeBuf I__1654 (
            .O(N__14167),
            .I(N__14161));
    CascadeBuf I__1653 (
            .O(N__14164),
            .I(N__14158));
    CascadeMux I__1652 (
            .O(N__14161),
            .I(N__14155));
    CascadeMux I__1651 (
            .O(N__14158),
            .I(N__14152));
    CascadeBuf I__1650 (
            .O(N__14155),
            .I(N__14149));
    CascadeBuf I__1649 (
            .O(N__14152),
            .I(N__14146));
    CascadeMux I__1648 (
            .O(N__14149),
            .I(N__14143));
    CascadeMux I__1647 (
            .O(N__14146),
            .I(N__14140));
    CascadeBuf I__1646 (
            .O(N__14143),
            .I(N__14137));
    InMux I__1645 (
            .O(N__14140),
            .I(N__14134));
    CascadeMux I__1644 (
            .O(N__14137),
            .I(N__14131));
    LocalMux I__1643 (
            .O(N__14134),
            .I(N__14128));
    InMux I__1642 (
            .O(N__14131),
            .I(N__14125));
    Span4Mux_s1_v I__1641 (
            .O(N__14128),
            .I(N__14116));
    LocalMux I__1640 (
            .O(N__14125),
            .I(N__14116));
    InMux I__1639 (
            .O(N__14124),
            .I(N__14113));
    CascadeMux I__1638 (
            .O(N__14123),
            .I(N__14110));
    CascadeMux I__1637 (
            .O(N__14122),
            .I(N__14107));
    CascadeMux I__1636 (
            .O(N__14121),
            .I(N__14104));
    Span4Mux_h I__1635 (
            .O(N__14116),
            .I(N__14101));
    LocalMux I__1634 (
            .O(N__14113),
            .I(N__14098));
    InMux I__1633 (
            .O(N__14110),
            .I(N__14095));
    InMux I__1632 (
            .O(N__14107),
            .I(N__14092));
    InMux I__1631 (
            .O(N__14104),
            .I(N__14089));
    Span4Mux_h I__1630 (
            .O(N__14101),
            .I(N__14086));
    Odrv4 I__1629 (
            .O(N__14098),
            .I(address_7));
    LocalMux I__1628 (
            .O(N__14095),
            .I(address_7));
    LocalMux I__1627 (
            .O(N__14092),
            .I(address_7));
    LocalMux I__1626 (
            .O(N__14089),
            .I(address_7));
    Odrv4 I__1625 (
            .O(N__14086),
            .I(address_7));
    InMux I__1624 (
            .O(N__14075),
            .I(N__14069));
    InMux I__1623 (
            .O(N__14074),
            .I(N__14069));
    LocalMux I__1622 (
            .O(N__14069),
            .I(N__14066));
    Odrv4 I__1621 (
            .O(N__14066),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_5 ));
    CascadeMux I__1620 (
            .O(N__14063),
            .I(N__14060));
    InMux I__1619 (
            .O(N__14060),
            .I(N__14054));
    InMux I__1618 (
            .O(N__14059),
            .I(N__14054));
    LocalMux I__1617 (
            .O(N__14054),
            .I(N__14051));
    Odrv4 I__1616 (
            .O(N__14051),
            .I(\processor_zipi8.pc_vector_5 ));
    InMux I__1615 (
            .O(N__14048),
            .I(N__14045));
    LocalMux I__1614 (
            .O(N__14045),
            .I(\processor_zipi8.program_counter_i.carry_pc_28_4 ));
    CascadeMux I__1613 (
            .O(N__14042),
            .I(N__14039));
    CascadeBuf I__1612 (
            .O(N__14039),
            .I(N__14035));
    CascadeMux I__1611 (
            .O(N__14038),
            .I(N__14032));
    CascadeMux I__1610 (
            .O(N__14035),
            .I(N__14029));
    CascadeBuf I__1609 (
            .O(N__14032),
            .I(N__14026));
    CascadeBuf I__1608 (
            .O(N__14029),
            .I(N__14023));
    CascadeMux I__1607 (
            .O(N__14026),
            .I(N__14020));
    CascadeMux I__1606 (
            .O(N__14023),
            .I(N__14017));
    CascadeBuf I__1605 (
            .O(N__14020),
            .I(N__14014));
    CascadeBuf I__1604 (
            .O(N__14017),
            .I(N__14011));
    CascadeMux I__1603 (
            .O(N__14014),
            .I(N__14008));
    CascadeMux I__1602 (
            .O(N__14011),
            .I(N__14005));
    CascadeBuf I__1601 (
            .O(N__14008),
            .I(N__14002));
    CascadeBuf I__1600 (
            .O(N__14005),
            .I(N__13999));
    CascadeMux I__1599 (
            .O(N__14002),
            .I(N__13996));
    CascadeMux I__1598 (
            .O(N__13999),
            .I(N__13993));
    CascadeBuf I__1597 (
            .O(N__13996),
            .I(N__13990));
    CascadeBuf I__1596 (
            .O(N__13993),
            .I(N__13987));
    CascadeMux I__1595 (
            .O(N__13990),
            .I(N__13984));
    CascadeMux I__1594 (
            .O(N__13987),
            .I(N__13981));
    CascadeBuf I__1593 (
            .O(N__13984),
            .I(N__13978));
    CascadeBuf I__1592 (
            .O(N__13981),
            .I(N__13975));
    CascadeMux I__1591 (
            .O(N__13978),
            .I(N__13972));
    CascadeMux I__1590 (
            .O(N__13975),
            .I(N__13969));
    CascadeBuf I__1589 (
            .O(N__13972),
            .I(N__13966));
    CascadeBuf I__1588 (
            .O(N__13969),
            .I(N__13963));
    CascadeMux I__1587 (
            .O(N__13966),
            .I(N__13960));
    CascadeMux I__1586 (
            .O(N__13963),
            .I(N__13957));
    CascadeBuf I__1585 (
            .O(N__13960),
            .I(N__13954));
    InMux I__1584 (
            .O(N__13957),
            .I(N__13951));
    CascadeMux I__1583 (
            .O(N__13954),
            .I(N__13948));
    LocalMux I__1582 (
            .O(N__13951),
            .I(N__13945));
    InMux I__1581 (
            .O(N__13948),
            .I(N__13942));
    Span4Mux_s1_v I__1580 (
            .O(N__13945),
            .I(N__13933));
    LocalMux I__1579 (
            .O(N__13942),
            .I(N__13933));
    InMux I__1578 (
            .O(N__13941),
            .I(N__13930));
    CascadeMux I__1577 (
            .O(N__13940),
            .I(N__13927));
    CascadeMux I__1576 (
            .O(N__13939),
            .I(N__13924));
    CascadeMux I__1575 (
            .O(N__13938),
            .I(N__13921));
    Span4Mux_h I__1574 (
            .O(N__13933),
            .I(N__13918));
    LocalMux I__1573 (
            .O(N__13930),
            .I(N__13915));
    InMux I__1572 (
            .O(N__13927),
            .I(N__13912));
    InMux I__1571 (
            .O(N__13924),
            .I(N__13909));
    InMux I__1570 (
            .O(N__13921),
            .I(N__13906));
    Span4Mux_h I__1569 (
            .O(N__13918),
            .I(N__13903));
    Odrv4 I__1568 (
            .O(N__13915),
            .I(address_5));
    LocalMux I__1567 (
            .O(N__13912),
            .I(address_5));
    LocalMux I__1566 (
            .O(N__13909),
            .I(address_5));
    LocalMux I__1565 (
            .O(N__13906),
            .I(address_5));
    Odrv4 I__1564 (
            .O(N__13903),
            .I(address_5));
    InMux I__1563 (
            .O(N__13892),
            .I(N__13889));
    LocalMux I__1562 (
            .O(N__13889),
            .I(N__13886));
    Odrv4 I__1561 (
            .O(N__13886),
            .I(\processor_zipi8.return_vector_11 ));
    CascadeMux I__1560 (
            .O(N__13883),
            .I(\processor_zipi8.program_counter_i.un3_half_pcZ0_cascade_ ));
    InMux I__1559 (
            .O(N__13880),
            .I(N__13874));
    InMux I__1558 (
            .O(N__13879),
            .I(N__13874));
    LocalMux I__1557 (
            .O(N__13874),
            .I(\processor_zipi8.flags_i.N_37 ));
    InMux I__1556 (
            .O(N__13871),
            .I(N__13868));
    LocalMux I__1555 (
            .O(N__13868),
            .I(\processor_zipi8.stack_memory_7 ));
    InMux I__1554 (
            .O(N__13865),
            .I(N__13862));
    LocalMux I__1553 (
            .O(N__13862),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_7 ));
    InMux I__1552 (
            .O(N__13859),
            .I(N__13856));
    LocalMux I__1551 (
            .O(N__13856),
            .I(N__13853));
    Span4Mux_v I__1550 (
            .O(N__13853),
            .I(N__13850));
    Odrv4 I__1549 (
            .O(N__13850),
            .I(\processor_zipi8.stack_memory_1 ));
    InMux I__1548 (
            .O(N__13847),
            .I(N__13844));
    LocalMux I__1547 (
            .O(N__13844),
            .I(N__13841));
    Span4Mux_v I__1546 (
            .O(N__13841),
            .I(N__13838));
    Odrv4 I__1545 (
            .O(N__13838),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_155 ));
    CascadeMux I__1544 (
            .O(N__13835),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_195_cascade_ ));
    CascadeMux I__1543 (
            .O(N__13832),
            .I(N__13828));
    CascadeMux I__1542 (
            .O(N__13831),
            .I(N__13825));
    CascadeBuf I__1541 (
            .O(N__13828),
            .I(N__13822));
    CascadeBuf I__1540 (
            .O(N__13825),
            .I(N__13819));
    CascadeMux I__1539 (
            .O(N__13822),
            .I(N__13816));
    CascadeMux I__1538 (
            .O(N__13819),
            .I(N__13813));
    CascadeBuf I__1537 (
            .O(N__13816),
            .I(N__13810));
    CascadeBuf I__1536 (
            .O(N__13813),
            .I(N__13807));
    CascadeMux I__1535 (
            .O(N__13810),
            .I(N__13804));
    CascadeMux I__1534 (
            .O(N__13807),
            .I(N__13801));
    CascadeBuf I__1533 (
            .O(N__13804),
            .I(N__13798));
    CascadeBuf I__1532 (
            .O(N__13801),
            .I(N__13795));
    CascadeMux I__1531 (
            .O(N__13798),
            .I(N__13792));
    CascadeMux I__1530 (
            .O(N__13795),
            .I(N__13789));
    CascadeBuf I__1529 (
            .O(N__13792),
            .I(N__13786));
    CascadeBuf I__1528 (
            .O(N__13789),
            .I(N__13783));
    CascadeMux I__1527 (
            .O(N__13786),
            .I(N__13780));
    CascadeMux I__1526 (
            .O(N__13783),
            .I(N__13777));
    CascadeBuf I__1525 (
            .O(N__13780),
            .I(N__13774));
    CascadeBuf I__1524 (
            .O(N__13777),
            .I(N__13771));
    CascadeMux I__1523 (
            .O(N__13774),
            .I(N__13768));
    CascadeMux I__1522 (
            .O(N__13771),
            .I(N__13765));
    CascadeBuf I__1521 (
            .O(N__13768),
            .I(N__13762));
    CascadeBuf I__1520 (
            .O(N__13765),
            .I(N__13759));
    CascadeMux I__1519 (
            .O(N__13762),
            .I(N__13756));
    CascadeMux I__1518 (
            .O(N__13759),
            .I(N__13753));
    CascadeBuf I__1517 (
            .O(N__13756),
            .I(N__13750));
    CascadeBuf I__1516 (
            .O(N__13753),
            .I(N__13747));
    CascadeMux I__1515 (
            .O(N__13750),
            .I(N__13744));
    CascadeMux I__1514 (
            .O(N__13747),
            .I(N__13741));
    InMux I__1513 (
            .O(N__13744),
            .I(N__13737));
    InMux I__1512 (
            .O(N__13741),
            .I(N__13734));
    InMux I__1511 (
            .O(N__13740),
            .I(N__13731));
    LocalMux I__1510 (
            .O(N__13737),
            .I(N__13723));
    LocalMux I__1509 (
            .O(N__13734),
            .I(N__13723));
    LocalMux I__1508 (
            .O(N__13731),
            .I(N__13720));
    InMux I__1507 (
            .O(N__13730),
            .I(N__13717));
    CascadeMux I__1506 (
            .O(N__13729),
            .I(N__13714));
    CascadeMux I__1505 (
            .O(N__13728),
            .I(N__13711));
    Span4Mux_v I__1504 (
            .O(N__13723),
            .I(N__13708));
    Span4Mux_h I__1503 (
            .O(N__13720),
            .I(N__13705));
    LocalMux I__1502 (
            .O(N__13717),
            .I(N__13702));
    InMux I__1501 (
            .O(N__13714),
            .I(N__13699));
    InMux I__1500 (
            .O(N__13711),
            .I(N__13696));
    Sp12to4 I__1499 (
            .O(N__13708),
            .I(N__13693));
    Odrv4 I__1498 (
            .O(N__13705),
            .I(address_6));
    Odrv4 I__1497 (
            .O(N__13702),
            .I(address_6));
    LocalMux I__1496 (
            .O(N__13699),
            .I(address_6));
    LocalMux I__1495 (
            .O(N__13696),
            .I(address_6));
    Odrv12 I__1494 (
            .O(N__13693),
            .I(address_6));
    CascadeMux I__1493 (
            .O(N__13682),
            .I(N__13678));
    CascadeMux I__1492 (
            .O(N__13681),
            .I(N__13675));
    CascadeBuf I__1491 (
            .O(N__13678),
            .I(N__13672));
    CascadeBuf I__1490 (
            .O(N__13675),
            .I(N__13669));
    CascadeMux I__1489 (
            .O(N__13672),
            .I(N__13666));
    CascadeMux I__1488 (
            .O(N__13669),
            .I(N__13663));
    CascadeBuf I__1487 (
            .O(N__13666),
            .I(N__13660));
    CascadeBuf I__1486 (
            .O(N__13663),
            .I(N__13657));
    CascadeMux I__1485 (
            .O(N__13660),
            .I(N__13654));
    CascadeMux I__1484 (
            .O(N__13657),
            .I(N__13651));
    CascadeBuf I__1483 (
            .O(N__13654),
            .I(N__13648));
    CascadeBuf I__1482 (
            .O(N__13651),
            .I(N__13645));
    CascadeMux I__1481 (
            .O(N__13648),
            .I(N__13642));
    CascadeMux I__1480 (
            .O(N__13645),
            .I(N__13639));
    CascadeBuf I__1479 (
            .O(N__13642),
            .I(N__13636));
    CascadeBuf I__1478 (
            .O(N__13639),
            .I(N__13633));
    CascadeMux I__1477 (
            .O(N__13636),
            .I(N__13630));
    CascadeMux I__1476 (
            .O(N__13633),
            .I(N__13627));
    CascadeBuf I__1475 (
            .O(N__13630),
            .I(N__13624));
    CascadeBuf I__1474 (
            .O(N__13627),
            .I(N__13621));
    CascadeMux I__1473 (
            .O(N__13624),
            .I(N__13618));
    CascadeMux I__1472 (
            .O(N__13621),
            .I(N__13615));
    CascadeBuf I__1471 (
            .O(N__13618),
            .I(N__13612));
    CascadeBuf I__1470 (
            .O(N__13615),
            .I(N__13609));
    CascadeMux I__1469 (
            .O(N__13612),
            .I(N__13606));
    CascadeMux I__1468 (
            .O(N__13609),
            .I(N__13603));
    CascadeBuf I__1467 (
            .O(N__13606),
            .I(N__13600));
    CascadeBuf I__1466 (
            .O(N__13603),
            .I(N__13597));
    CascadeMux I__1465 (
            .O(N__13600),
            .I(N__13593));
    CascadeMux I__1464 (
            .O(N__13597),
            .I(N__13590));
    InMux I__1463 (
            .O(N__13596),
            .I(N__13587));
    InMux I__1462 (
            .O(N__13593),
            .I(N__13581));
    InMux I__1461 (
            .O(N__13590),
            .I(N__13578));
    LocalMux I__1460 (
            .O(N__13587),
            .I(N__13575));
    CascadeMux I__1459 (
            .O(N__13586),
            .I(N__13572));
    CascadeMux I__1458 (
            .O(N__13585),
            .I(N__13569));
    CascadeMux I__1457 (
            .O(N__13584),
            .I(N__13566));
    LocalMux I__1456 (
            .O(N__13581),
            .I(N__13561));
    LocalMux I__1455 (
            .O(N__13578),
            .I(N__13561));
    Span4Mux_h I__1454 (
            .O(N__13575),
            .I(N__13558));
    InMux I__1453 (
            .O(N__13572),
            .I(N__13555));
    InMux I__1452 (
            .O(N__13569),
            .I(N__13552));
    InMux I__1451 (
            .O(N__13566),
            .I(N__13549));
    Span12Mux_s4_v I__1450 (
            .O(N__13561),
            .I(N__13546));
    Odrv4 I__1449 (
            .O(N__13558),
            .I(address_4));
    LocalMux I__1448 (
            .O(N__13555),
            .I(address_4));
    LocalMux I__1447 (
            .O(N__13552),
            .I(address_4));
    LocalMux I__1446 (
            .O(N__13549),
            .I(address_4));
    Odrv12 I__1445 (
            .O(N__13546),
            .I(address_4));
    InMux I__1444 (
            .O(N__13535),
            .I(N__13532));
    LocalMux I__1443 (
            .O(N__13532),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_4 ));
    InMux I__1442 (
            .O(N__13529),
            .I(N__13526));
    LocalMux I__1441 (
            .O(N__13526),
            .I(N__13523));
    Odrv4 I__1440 (
            .O(N__13523),
            .I(\processor_zipi8.stack_memory_6 ));
    InMux I__1439 (
            .O(N__13520),
            .I(N__13517));
    LocalMux I__1438 (
            .O(N__13517),
            .I(N__13514));
    Odrv4 I__1437 (
            .O(N__13514),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_6 ));
    CascadeMux I__1436 (
            .O(N__13511),
            .I(\processor_zipi8.flags_i.N_125_mux_cascade_ ));
    InMux I__1435 (
            .O(N__13508),
            .I(N__13505));
    LocalMux I__1434 (
            .O(N__13505),
            .I(\processor_zipi8.stack_i.stack_bit ));
    InMux I__1433 (
            .O(N__13502),
            .I(N__13497));
    InMux I__1432 (
            .O(N__13501),
            .I(N__13492));
    InMux I__1431 (
            .O(N__13500),
            .I(N__13492));
    LocalMux I__1430 (
            .O(N__13497),
            .I(\processor_zipi8.run ));
    LocalMux I__1429 (
            .O(N__13492),
            .I(\processor_zipi8.run ));
    InMux I__1428 (
            .O(N__13487),
            .I(N__13481));
    InMux I__1427 (
            .O(N__13486),
            .I(N__13481));
    LocalMux I__1426 (
            .O(N__13481),
            .I(N__13478));
    Span4Mux_v I__1425 (
            .O(N__13478),
            .I(N__13475));
    Span4Mux_h I__1424 (
            .O(N__13475),
            .I(N__13472));
    Span4Mux_h I__1423 (
            .O(N__13472),
            .I(N__13469));
    Odrv4 I__1422 (
            .O(N__13469),
            .I(BTN1_c));
    InMux I__1421 (
            .O(N__13466),
            .I(N__13463));
    LocalMux I__1420 (
            .O(N__13463),
            .I(\processor_zipi8.stack_memory_2 ));
    CascadeMux I__1419 (
            .O(N__13460),
            .I(N__13456));
    InMux I__1418 (
            .O(N__13459),
            .I(N__13451));
    InMux I__1417 (
            .O(N__13456),
            .I(N__13451));
    LocalMux I__1416 (
            .O(N__13451),
            .I(\processor_zipi8.special_bit ));
    IoInMux I__1415 (
            .O(N__13448),
            .I(N__13445));
    LocalMux I__1414 (
            .O(N__13445),
            .I(N__13442));
    Span4Mux_s1_h I__1413 (
            .O(N__13442),
            .I(N__13439));
    Odrv4 I__1412 (
            .O(N__13439),
            .I(\processor_zipi8.state_machine_i.bram_enable ));
    InMux I__1411 (
            .O(N__13436),
            .I(N__13433));
    LocalMux I__1410 (
            .O(N__13433),
            .I(\processor_zipi8.stack_memory_11 ));
    InMux I__1409 (
            .O(N__13430),
            .I(N__13424));
    InMux I__1408 (
            .O(N__13429),
            .I(N__13424));
    LocalMux I__1407 (
            .O(N__13424),
            .I(N__13421));
    Span4Mux_v I__1406 (
            .O(N__13421),
            .I(N__13418));
    Odrv4 I__1405 (
            .O(N__13418),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_6 ));
    CascadeMux I__1404 (
            .O(N__13415),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_6_cascade_ ));
    InMux I__1403 (
            .O(N__13412),
            .I(N__13409));
    LocalMux I__1402 (
            .O(N__13409),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_6 ));
    InMux I__1401 (
            .O(N__13406),
            .I(N__13402));
    InMux I__1400 (
            .O(N__13405),
            .I(N__13399));
    LocalMux I__1399 (
            .O(N__13402),
            .I(N__13396));
    LocalMux I__1398 (
            .O(N__13399),
            .I(N__13393));
    Span4Mux_v I__1397 (
            .O(N__13396),
            .I(N__13390));
    Span4Mux_v I__1396 (
            .O(N__13393),
            .I(N__13387));
    Span4Mux_v I__1395 (
            .O(N__13390),
            .I(N__13384));
    Odrv4 I__1394 (
            .O(N__13387),
            .I(\processor_zipi8.sy_6 ));
    Odrv4 I__1393 (
            .O(N__13384),
            .I(\processor_zipi8.sy_6 ));
    CascadeMux I__1392 (
            .O(N__13379),
            .I(\processor_zipi8.port_id_6_cascade_ ));
    InMux I__1391 (
            .O(N__13376),
            .I(N__13373));
    LocalMux I__1390 (
            .O(N__13373),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_6 ));
    CascadeMux I__1389 (
            .O(N__13370),
            .I(N__13367));
    InMux I__1388 (
            .O(N__13367),
            .I(N__13363));
    CascadeMux I__1387 (
            .O(N__13366),
            .I(N__13359));
    LocalMux I__1386 (
            .O(N__13363),
            .I(N__13356));
    CascadeMux I__1385 (
            .O(N__13362),
            .I(N__13352));
    InMux I__1384 (
            .O(N__13359),
            .I(N__13348));
    Span4Mux_v I__1383 (
            .O(N__13356),
            .I(N__13345));
    InMux I__1382 (
            .O(N__13355),
            .I(N__13338));
    InMux I__1381 (
            .O(N__13352),
            .I(N__13338));
    InMux I__1380 (
            .O(N__13351),
            .I(N__13338));
    LocalMux I__1379 (
            .O(N__13348),
            .I(\processor_zipi8.port_id_6 ));
    Odrv4 I__1378 (
            .O(N__13345),
            .I(\processor_zipi8.port_id_6 ));
    LocalMux I__1377 (
            .O(N__13338),
            .I(\processor_zipi8.port_id_6 ));
    InMux I__1376 (
            .O(N__13331),
            .I(N__13328));
    LocalMux I__1375 (
            .O(N__13328),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_6 ));
    InMux I__1374 (
            .O(N__13325),
            .I(N__13319));
    InMux I__1373 (
            .O(N__13324),
            .I(N__13319));
    LocalMux I__1372 (
            .O(N__13319),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_5 ));
    InMux I__1371 (
            .O(N__13316),
            .I(N__13312));
    InMux I__1370 (
            .O(N__13315),
            .I(N__13309));
    LocalMux I__1369 (
            .O(N__13312),
            .I(N__13304));
    LocalMux I__1368 (
            .O(N__13309),
            .I(N__13304));
    Odrv12 I__1367 (
            .O(N__13304),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_6 ));
    InMux I__1366 (
            .O(N__13301),
            .I(N__13295));
    InMux I__1365 (
            .O(N__13300),
            .I(N__13295));
    LocalMux I__1364 (
            .O(N__13295),
            .I(N__13292));
    Odrv4 I__1363 (
            .O(N__13292),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_7 ));
    InMux I__1362 (
            .O(N__13289),
            .I(N__13286));
    LocalMux I__1361 (
            .O(N__13286),
            .I(\processor_zipi8.spm_data_5 ));
    CascadeMux I__1360 (
            .O(N__13283),
            .I(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202_cascade_ ));
    InMux I__1359 (
            .O(N__13280),
            .I(N__13274));
    InMux I__1358 (
            .O(N__13279),
            .I(N__13274));
    LocalMux I__1357 (
            .O(N__13274),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_5 ));
    CascadeMux I__1356 (
            .O(N__13271),
            .I(N__13268));
    InMux I__1355 (
            .O(N__13268),
            .I(N__13265));
    LocalMux I__1354 (
            .O(N__13265),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_5 ));
    InMux I__1353 (
            .O(N__13262),
            .I(N__13256));
    InMux I__1352 (
            .O(N__13261),
            .I(N__13256));
    LocalMux I__1351 (
            .O(N__13256),
            .I(N__13253));
    Odrv4 I__1350 (
            .O(N__13253),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_6 ));
    InMux I__1349 (
            .O(N__13250),
            .I(N__13247));
    LocalMux I__1348 (
            .O(N__13247),
            .I(N__13244));
    Span4Mux_s2_h I__1347 (
            .O(N__13244),
            .I(N__13240));
    InMux I__1346 (
            .O(N__13243),
            .I(N__13237));
    Odrv4 I__1345 (
            .O(N__13240),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7 ));
    LocalMux I__1344 (
            .O(N__13237),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7 ));
    InMux I__1343 (
            .O(N__13232),
            .I(N__13229));
    LocalMux I__1342 (
            .O(N__13229),
            .I(N__13226));
    Odrv4 I__1341 (
            .O(N__13226),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_7 ));
    InMux I__1340 (
            .O(N__13223),
            .I(N__13217));
    InMux I__1339 (
            .O(N__13222),
            .I(N__13217));
    LocalMux I__1338 (
            .O(N__13217),
            .I(N__13214));
    Odrv4 I__1337 (
            .O(N__13214),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_5 ));
    InMux I__1336 (
            .O(N__13211),
            .I(N__13205));
    InMux I__1335 (
            .O(N__13210),
            .I(N__13205));
    LocalMux I__1334 (
            .O(N__13205),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_6 ));
    InMux I__1333 (
            .O(N__13202),
            .I(N__13198));
    InMux I__1332 (
            .O(N__13201),
            .I(N__13195));
    LocalMux I__1331 (
            .O(N__13198),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7 ));
    LocalMux I__1330 (
            .O(N__13195),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7 ));
    CascadeMux I__1329 (
            .O(N__13190),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_6_cascade_ ));
    InMux I__1328 (
            .O(N__13187),
            .I(N__13184));
    LocalMux I__1327 (
            .O(N__13184),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_6 ));
    CascadeMux I__1326 (
            .O(N__13181),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_6_cascade_ ));
    InMux I__1325 (
            .O(N__13178),
            .I(N__13175));
    LocalMux I__1324 (
            .O(N__13175),
            .I(N__13172));
    Odrv4 I__1323 (
            .O(N__13172),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_6 ));
    CascadeMux I__1322 (
            .O(N__13169),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_6_cascade_ ));
    InMux I__1321 (
            .O(N__13166),
            .I(N__13163));
    LocalMux I__1320 (
            .O(N__13163),
            .I(N__13160));
    Odrv4 I__1319 (
            .O(N__13160),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_6 ));
    CascadeMux I__1318 (
            .O(N__13157),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_6_cascade_ ));
    CascadeMux I__1317 (
            .O(N__13154),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_6_cascade_ ));
    InMux I__1316 (
            .O(N__13151),
            .I(N__13147));
    InMux I__1315 (
            .O(N__13150),
            .I(N__13144));
    LocalMux I__1314 (
            .O(N__13147),
            .I(N__13139));
    LocalMux I__1313 (
            .O(N__13144),
            .I(N__13139));
    Span4Mux_v I__1312 (
            .O(N__13139),
            .I(N__13136));
    Odrv4 I__1311 (
            .O(N__13136),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_7 ));
    CascadeMux I__1310 (
            .O(N__13133),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_6_cascade_ ));
    InMux I__1309 (
            .O(N__13130),
            .I(N__13126));
    InMux I__1308 (
            .O(N__13129),
            .I(N__13123));
    LocalMux I__1307 (
            .O(N__13126),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6 ));
    LocalMux I__1306 (
            .O(N__13123),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6 ));
    CascadeMux I__1305 (
            .O(N__13118),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_7_cascade_ ));
    InMux I__1304 (
            .O(N__13115),
            .I(N__13112));
    LocalMux I__1303 (
            .O(N__13112),
            .I(N__13109));
    Span4Mux_v I__1302 (
            .O(N__13109),
            .I(N__13106));
    Odrv4 I__1301 (
            .O(N__13106),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIK2TR1_7 ));
    InMux I__1300 (
            .O(N__13103),
            .I(N__13099));
    InMux I__1299 (
            .O(N__13102),
            .I(N__13096));
    LocalMux I__1298 (
            .O(N__13099),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7 ));
    LocalMux I__1297 (
            .O(N__13096),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7 ));
    InMux I__1296 (
            .O(N__13091),
            .I(N__13088));
    LocalMux I__1295 (
            .O(N__13088),
            .I(\processor_zipi8.alu_result_3 ));
    CascadeMux I__1294 (
            .O(N__13085),
            .I(\processor_zipi8.flags_i.m82_1_cascade_ ));
    InMux I__1293 (
            .O(N__13082),
            .I(N__13079));
    LocalMux I__1292 (
            .O(N__13079),
            .I(\processor_zipi8.flags_i.m82_1 ));
    CascadeMux I__1291 (
            .O(N__13076),
            .I(N__13073));
    InMux I__1290 (
            .O(N__13073),
            .I(N__13070));
    LocalMux I__1289 (
            .O(N__13070),
            .I(N__13067));
    Span4Mux_h I__1288 (
            .O(N__13067),
            .I(N__13064));
    Span4Mux_v I__1287 (
            .O(N__13064),
            .I(N__13061));
    Odrv4 I__1286 (
            .O(N__13061),
            .I(\processor_zipi8.zero_flag_RNIJSPM4 ));
    InMux I__1285 (
            .O(N__13058),
            .I(N__13055));
    LocalMux I__1284 (
            .O(N__13055),
            .I(\processor_zipi8.flags_i.N_55 ));
    CascadeMux I__1283 (
            .O(N__13052),
            .I(\processor_zipi8.flags_i.m61_ns_1_cascade_ ));
    InMux I__1282 (
            .O(N__13049),
            .I(N__13046));
    LocalMux I__1281 (
            .O(N__13046),
            .I(N__13043));
    Odrv4 I__1280 (
            .O(N__13043),
            .I(\processor_zipi8.pc_vector_8 ));
    CascadeMux I__1279 (
            .O(N__13040),
            .I(\processor_zipi8.program_counter_i.carry_pc_46_7_cascade_ ));
    CascadeMux I__1278 (
            .O(N__13037),
            .I(N__13033));
    CascadeMux I__1277 (
            .O(N__13036),
            .I(N__13030));
    CascadeBuf I__1276 (
            .O(N__13033),
            .I(N__13027));
    CascadeBuf I__1275 (
            .O(N__13030),
            .I(N__13024));
    CascadeMux I__1274 (
            .O(N__13027),
            .I(N__13021));
    CascadeMux I__1273 (
            .O(N__13024),
            .I(N__13018));
    CascadeBuf I__1272 (
            .O(N__13021),
            .I(N__13015));
    CascadeBuf I__1271 (
            .O(N__13018),
            .I(N__13012));
    CascadeMux I__1270 (
            .O(N__13015),
            .I(N__13009));
    CascadeMux I__1269 (
            .O(N__13012),
            .I(N__13006));
    CascadeBuf I__1268 (
            .O(N__13009),
            .I(N__13003));
    CascadeBuf I__1267 (
            .O(N__13006),
            .I(N__13000));
    CascadeMux I__1266 (
            .O(N__13003),
            .I(N__12997));
    CascadeMux I__1265 (
            .O(N__13000),
            .I(N__12994));
    CascadeBuf I__1264 (
            .O(N__12997),
            .I(N__12991));
    CascadeBuf I__1263 (
            .O(N__12994),
            .I(N__12988));
    CascadeMux I__1262 (
            .O(N__12991),
            .I(N__12985));
    CascadeMux I__1261 (
            .O(N__12988),
            .I(N__12982));
    CascadeBuf I__1260 (
            .O(N__12985),
            .I(N__12979));
    CascadeBuf I__1259 (
            .O(N__12982),
            .I(N__12976));
    CascadeMux I__1258 (
            .O(N__12979),
            .I(N__12973));
    CascadeMux I__1257 (
            .O(N__12976),
            .I(N__12970));
    CascadeBuf I__1256 (
            .O(N__12973),
            .I(N__12967));
    CascadeBuf I__1255 (
            .O(N__12970),
            .I(N__12964));
    CascadeMux I__1254 (
            .O(N__12967),
            .I(N__12961));
    CascadeMux I__1253 (
            .O(N__12964),
            .I(N__12958));
    CascadeBuf I__1252 (
            .O(N__12961),
            .I(N__12955));
    CascadeBuf I__1251 (
            .O(N__12958),
            .I(N__12952));
    CascadeMux I__1250 (
            .O(N__12955),
            .I(N__12948));
    CascadeMux I__1249 (
            .O(N__12952),
            .I(N__12945));
    CascadeMux I__1248 (
            .O(N__12951),
            .I(N__12940));
    InMux I__1247 (
            .O(N__12948),
            .I(N__12936));
    InMux I__1246 (
            .O(N__12945),
            .I(N__12933));
    InMux I__1245 (
            .O(N__12944),
            .I(N__12930));
    CascadeMux I__1244 (
            .O(N__12943),
            .I(N__12927));
    InMux I__1243 (
            .O(N__12940),
            .I(N__12924));
    CascadeMux I__1242 (
            .O(N__12939),
            .I(N__12921));
    LocalMux I__1241 (
            .O(N__12936),
            .I(N__12918));
    LocalMux I__1240 (
            .O(N__12933),
            .I(N__12915));
    LocalMux I__1239 (
            .O(N__12930),
            .I(N__12912));
    InMux I__1238 (
            .O(N__12927),
            .I(N__12909));
    LocalMux I__1237 (
            .O(N__12924),
            .I(N__12906));
    InMux I__1236 (
            .O(N__12921),
            .I(N__12903));
    Span4Mux_v I__1235 (
            .O(N__12918),
            .I(N__12898));
    Span4Mux_v I__1234 (
            .O(N__12915),
            .I(N__12898));
    Span4Mux_h I__1233 (
            .O(N__12912),
            .I(N__12895));
    LocalMux I__1232 (
            .O(N__12909),
            .I(N__12890));
    Span4Mux_h I__1231 (
            .O(N__12906),
            .I(N__12890));
    LocalMux I__1230 (
            .O(N__12903),
            .I(N__12885));
    Sp12to4 I__1229 (
            .O(N__12898),
            .I(N__12885));
    Odrv4 I__1228 (
            .O(N__12895),
            .I(address_8));
    Odrv4 I__1227 (
            .O(N__12890),
            .I(address_8));
    Odrv12 I__1226 (
            .O(N__12885),
            .I(address_8));
    InMux I__1225 (
            .O(N__12878),
            .I(N__12875));
    LocalMux I__1224 (
            .O(N__12875),
            .I(N__12871));
    InMux I__1223 (
            .O(N__12874),
            .I(N__12868));
    Odrv4 I__1222 (
            .O(N__12871),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_8 ));
    LocalMux I__1221 (
            .O(N__12868),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_8 ));
    CascadeMux I__1220 (
            .O(N__12863),
            .I(\processor_zipi8.flags_i.zero_flag_3_cascade_ ));
    CascadeMux I__1219 (
            .O(N__12860),
            .I(N__12857));
    InMux I__1218 (
            .O(N__12857),
            .I(N__12854));
    LocalMux I__1217 (
            .O(N__12854),
            .I(\processor_zipi8.shadow_zero_flag ));
    InMux I__1216 (
            .O(N__12851),
            .I(N__12848));
    LocalMux I__1215 (
            .O(N__12848),
            .I(N__12845));
    Span12Mux_s3_v I__1214 (
            .O(N__12845),
            .I(N__12842));
    Odrv12 I__1213 (
            .O(N__12842),
            .I(\processor_zipi8.alu_result_7 ));
    CascadeMux I__1212 (
            .O(N__12839),
            .I(\processor_zipi8.alu_result_6_cascade_ ));
    InMux I__1211 (
            .O(N__12836),
            .I(N__12833));
    LocalMux I__1210 (
            .O(N__12833),
            .I(\processor_zipi8.flags_i.zero_flag_3_0_5 ));
    InMux I__1209 (
            .O(N__12830),
            .I(N__12827));
    LocalMux I__1208 (
            .O(N__12827),
            .I(\processor_zipi8.alu_result_5 ));
    InMux I__1207 (
            .O(N__12824),
            .I(N__12821));
    LocalMux I__1206 (
            .O(N__12821),
            .I(N__12818));
    Span4Mux_s3_v I__1205 (
            .O(N__12818),
            .I(N__12815));
    Span4Mux_v I__1204 (
            .O(N__12815),
            .I(N__12812));
    Odrv4 I__1203 (
            .O(N__12812),
            .I(\processor_zipi8.stack_i.stack_zero_flag ));
    InMux I__1202 (
            .O(N__12809),
            .I(N__12806));
    LocalMux I__1201 (
            .O(N__12806),
            .I(\processor_zipi8.stack_i.shadow_zero_value ));
    InMux I__1200 (
            .O(N__12803),
            .I(N__12800));
    LocalMux I__1199 (
            .O(N__12800),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_8 ));
    CascadeMux I__1198 (
            .O(N__12797),
            .I(\processor_zipi8.pc_vector_8_cascade_ ));
    CascadeMux I__1197 (
            .O(N__12794),
            .I(\processor_zipi8.program_counter_i.half_pc_0_0_9_cascade_ ));
    CascadeMux I__1196 (
            .O(N__12791),
            .I(N__12787));
    CascadeMux I__1195 (
            .O(N__12790),
            .I(N__12784));
    CascadeBuf I__1194 (
            .O(N__12787),
            .I(N__12781));
    CascadeBuf I__1193 (
            .O(N__12784),
            .I(N__12778));
    CascadeMux I__1192 (
            .O(N__12781),
            .I(N__12775));
    CascadeMux I__1191 (
            .O(N__12778),
            .I(N__12772));
    CascadeBuf I__1190 (
            .O(N__12775),
            .I(N__12769));
    CascadeBuf I__1189 (
            .O(N__12772),
            .I(N__12766));
    CascadeMux I__1188 (
            .O(N__12769),
            .I(N__12763));
    CascadeMux I__1187 (
            .O(N__12766),
            .I(N__12760));
    CascadeBuf I__1186 (
            .O(N__12763),
            .I(N__12757));
    CascadeBuf I__1185 (
            .O(N__12760),
            .I(N__12754));
    CascadeMux I__1184 (
            .O(N__12757),
            .I(N__12751));
    CascadeMux I__1183 (
            .O(N__12754),
            .I(N__12748));
    CascadeBuf I__1182 (
            .O(N__12751),
            .I(N__12745));
    CascadeBuf I__1181 (
            .O(N__12748),
            .I(N__12742));
    CascadeMux I__1180 (
            .O(N__12745),
            .I(N__12739));
    CascadeMux I__1179 (
            .O(N__12742),
            .I(N__12736));
    CascadeBuf I__1178 (
            .O(N__12739),
            .I(N__12733));
    CascadeBuf I__1177 (
            .O(N__12736),
            .I(N__12730));
    CascadeMux I__1176 (
            .O(N__12733),
            .I(N__12727));
    CascadeMux I__1175 (
            .O(N__12730),
            .I(N__12724));
    CascadeBuf I__1174 (
            .O(N__12727),
            .I(N__12721));
    CascadeBuf I__1173 (
            .O(N__12724),
            .I(N__12718));
    CascadeMux I__1172 (
            .O(N__12721),
            .I(N__12715));
    CascadeMux I__1171 (
            .O(N__12718),
            .I(N__12712));
    CascadeBuf I__1170 (
            .O(N__12715),
            .I(N__12709));
    CascadeBuf I__1169 (
            .O(N__12712),
            .I(N__12706));
    CascadeMux I__1168 (
            .O(N__12709),
            .I(N__12703));
    CascadeMux I__1167 (
            .O(N__12706),
            .I(N__12700));
    InMux I__1166 (
            .O(N__12703),
            .I(N__12696));
    InMux I__1165 (
            .O(N__12700),
            .I(N__12693));
    CascadeMux I__1164 (
            .O(N__12699),
            .I(N__12688));
    LocalMux I__1163 (
            .O(N__12696),
            .I(N__12685));
    LocalMux I__1162 (
            .O(N__12693),
            .I(N__12682));
    InMux I__1161 (
            .O(N__12692),
            .I(N__12679));
    CascadeMux I__1160 (
            .O(N__12691),
            .I(N__12675));
    InMux I__1159 (
            .O(N__12688),
            .I(N__12672));
    Span4Mux_s1_v I__1158 (
            .O(N__12685),
            .I(N__12667));
    Span4Mux_s2_h I__1157 (
            .O(N__12682),
            .I(N__12667));
    LocalMux I__1156 (
            .O(N__12679),
            .I(N__12664));
    InMux I__1155 (
            .O(N__12678),
            .I(N__12661));
    InMux I__1154 (
            .O(N__12675),
            .I(N__12658));
    LocalMux I__1153 (
            .O(N__12672),
            .I(N__12655));
    Span4Mux_h I__1152 (
            .O(N__12667),
            .I(N__12652));
    Span4Mux_v I__1151 (
            .O(N__12664),
            .I(N__12645));
    LocalMux I__1150 (
            .O(N__12661),
            .I(N__12645));
    LocalMux I__1149 (
            .O(N__12658),
            .I(N__12645));
    Span4Mux_h I__1148 (
            .O(N__12655),
            .I(N__12640));
    Span4Mux_h I__1147 (
            .O(N__12652),
            .I(N__12640));
    Odrv4 I__1146 (
            .O(N__12645),
            .I(address_9));
    Odrv4 I__1145 (
            .O(N__12640),
            .I(address_9));
    CascadeMux I__1144 (
            .O(N__12635),
            .I(\processor_zipi8.program_counter_i.un380_half_pc_cascade_ ));
    CascadeMux I__1143 (
            .O(N__12632),
            .I(\processor_zipi8.program_counter_i.half_pc_0_10_cascade_ ));
    CascadeMux I__1142 (
            .O(N__12629),
            .I(N__12625));
    CascadeMux I__1141 (
            .O(N__12628),
            .I(N__12622));
    CascadeBuf I__1140 (
            .O(N__12625),
            .I(N__12619));
    CascadeBuf I__1139 (
            .O(N__12622),
            .I(N__12616));
    CascadeMux I__1138 (
            .O(N__12619),
            .I(N__12613));
    CascadeMux I__1137 (
            .O(N__12616),
            .I(N__12610));
    CascadeBuf I__1136 (
            .O(N__12613),
            .I(N__12607));
    CascadeBuf I__1135 (
            .O(N__12610),
            .I(N__12604));
    CascadeMux I__1134 (
            .O(N__12607),
            .I(N__12601));
    CascadeMux I__1133 (
            .O(N__12604),
            .I(N__12598));
    CascadeBuf I__1132 (
            .O(N__12601),
            .I(N__12595));
    CascadeBuf I__1131 (
            .O(N__12598),
            .I(N__12592));
    CascadeMux I__1130 (
            .O(N__12595),
            .I(N__12589));
    CascadeMux I__1129 (
            .O(N__12592),
            .I(N__12586));
    CascadeBuf I__1128 (
            .O(N__12589),
            .I(N__12583));
    CascadeBuf I__1127 (
            .O(N__12586),
            .I(N__12580));
    CascadeMux I__1126 (
            .O(N__12583),
            .I(N__12577));
    CascadeMux I__1125 (
            .O(N__12580),
            .I(N__12574));
    CascadeBuf I__1124 (
            .O(N__12577),
            .I(N__12571));
    CascadeBuf I__1123 (
            .O(N__12574),
            .I(N__12568));
    CascadeMux I__1122 (
            .O(N__12571),
            .I(N__12565));
    CascadeMux I__1121 (
            .O(N__12568),
            .I(N__12562));
    CascadeBuf I__1120 (
            .O(N__12565),
            .I(N__12559));
    CascadeBuf I__1119 (
            .O(N__12562),
            .I(N__12556));
    CascadeMux I__1118 (
            .O(N__12559),
            .I(N__12553));
    CascadeMux I__1117 (
            .O(N__12556),
            .I(N__12550));
    CascadeBuf I__1116 (
            .O(N__12553),
            .I(N__12547));
    CascadeBuf I__1115 (
            .O(N__12550),
            .I(N__12544));
    CascadeMux I__1114 (
            .O(N__12547),
            .I(N__12540));
    CascadeMux I__1113 (
            .O(N__12544),
            .I(N__12537));
    InMux I__1112 (
            .O(N__12543),
            .I(N__12533));
    InMux I__1111 (
            .O(N__12540),
            .I(N__12529));
    InMux I__1110 (
            .O(N__12537),
            .I(N__12526));
    CascadeMux I__1109 (
            .O(N__12536),
            .I(N__12523));
    LocalMux I__1108 (
            .O(N__12533),
            .I(N__12520));
    CascadeMux I__1107 (
            .O(N__12532),
            .I(N__12517));
    LocalMux I__1106 (
            .O(N__12529),
            .I(N__12512));
    LocalMux I__1105 (
            .O(N__12526),
            .I(N__12512));
    InMux I__1104 (
            .O(N__12523),
            .I(N__12509));
    Span4Mux_v I__1103 (
            .O(N__12520),
            .I(N__12506));
    InMux I__1102 (
            .O(N__12517),
            .I(N__12503));
    Span4Mux_s3_v I__1101 (
            .O(N__12512),
            .I(N__12500));
    LocalMux I__1100 (
            .O(N__12509),
            .I(N__12495));
    Sp12to4 I__1099 (
            .O(N__12506),
            .I(N__12490));
    LocalMux I__1098 (
            .O(N__12503),
            .I(N__12490));
    Span4Mux_h I__1097 (
            .O(N__12500),
            .I(N__12487));
    InMux I__1096 (
            .O(N__12499),
            .I(N__12482));
    InMux I__1095 (
            .O(N__12498),
            .I(N__12482));
    Span4Mux_h I__1094 (
            .O(N__12495),
            .I(N__12479));
    Span12Mux_s11_h I__1093 (
            .O(N__12490),
            .I(N__12476));
    Span4Mux_h I__1092 (
            .O(N__12487),
            .I(N__12473));
    LocalMux I__1091 (
            .O(N__12482),
            .I(address_10));
    Odrv4 I__1090 (
            .O(N__12479),
            .I(address_10));
    Odrv12 I__1089 (
            .O(N__12476),
            .I(address_10));
    Odrv4 I__1088 (
            .O(N__12473),
            .I(address_10));
    CascadeMux I__1087 (
            .O(N__12464),
            .I(N__12461));
    InMux I__1086 (
            .O(N__12461),
            .I(N__12458));
    LocalMux I__1085 (
            .O(N__12458),
            .I(N__12455));
    Span4Mux_v I__1084 (
            .O(N__12455),
            .I(N__12452));
    Odrv4 I__1083 (
            .O(N__12452),
            .I(\processor_zipi8.return_vector_10 ));
    InMux I__1082 (
            .O(N__12449),
            .I(N__12446));
    LocalMux I__1081 (
            .O(N__12446),
            .I(\processor_zipi8.program_counter_i.un395_half_pcZ0 ));
    InMux I__1080 (
            .O(N__12443),
            .I(N__12440));
    LocalMux I__1079 (
            .O(N__12440),
            .I(\processor_zipi8.program_counter_i.carry_pc_46_7 ));
    InMux I__1078 (
            .O(N__12437),
            .I(N__12434));
    LocalMux I__1077 (
            .O(N__12434),
            .I(N__12431));
    Odrv4 I__1076 (
            .O(N__12431),
            .I(\processor_zipi8.stack_memory_9 ));
    InMux I__1075 (
            .O(N__12428),
            .I(N__12425));
    LocalMux I__1074 (
            .O(N__12425),
            .I(N__12422));
    Odrv4 I__1073 (
            .O(N__12422),
            .I(\processor_zipi8.stack_memory_4 ));
    InMux I__1072 (
            .O(N__12419),
            .I(N__12416));
    LocalMux I__1071 (
            .O(N__12416),
            .I(N__12413));
    Span4Mux_v I__1070 (
            .O(N__12413),
            .I(N__12410));
    Odrv4 I__1069 (
            .O(N__12410),
            .I(\processor_zipi8.stack_memory_8 ));
    InMux I__1068 (
            .O(N__12407),
            .I(N__12404));
    LocalMux I__1067 (
            .O(N__12404),
            .I(N__12401));
    Span4Mux_v I__1066 (
            .O(N__12401),
            .I(N__12398));
    Odrv4 I__1065 (
            .O(N__12398),
            .I(\processor_zipi8.stack_memory_10 ));
    InMux I__1064 (
            .O(N__12395),
            .I(N__12392));
    LocalMux I__1063 (
            .O(N__12392),
            .I(N__12389));
    Span4Mux_h I__1062 (
            .O(N__12389),
            .I(N__12386));
    Odrv4 I__1061 (
            .O(N__12386),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_9 ));
    InMux I__1060 (
            .O(N__12383),
            .I(N__12379));
    InMux I__1059 (
            .O(N__12382),
            .I(N__12376));
    LocalMux I__1058 (
            .O(N__12379),
            .I(N__12371));
    LocalMux I__1057 (
            .O(N__12376),
            .I(N__12371));
    Odrv12 I__1056 (
            .O(N__12371),
            .I(\processor_zipi8.sy_5 ));
    InMux I__1055 (
            .O(N__12368),
            .I(N__12364));
    InMux I__1054 (
            .O(N__12367),
            .I(N__12361));
    LocalMux I__1053 (
            .O(N__12364),
            .I(N__12358));
    LocalMux I__1052 (
            .O(N__12361),
            .I(N__12355));
    Span4Mux_h I__1051 (
            .O(N__12358),
            .I(N__12350));
    Span4Mux_v I__1050 (
            .O(N__12355),
            .I(N__12350));
    Odrv4 I__1049 (
            .O(N__12350),
            .I(\processor_zipi8.sy_7 ));
    InMux I__1048 (
            .O(N__12347),
            .I(N__12344));
    LocalMux I__1047 (
            .O(N__12344),
            .I(N__12341));
    Odrv4 I__1046 (
            .O(N__12341),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_7 ));
    InMux I__1045 (
            .O(N__12338),
            .I(N__12335));
    LocalMux I__1044 (
            .O(N__12335),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_7 ));
    CascadeMux I__1043 (
            .O(N__12332),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_7_cascade_ ));
    InMux I__1042 (
            .O(N__12329),
            .I(N__12326));
    LocalMux I__1041 (
            .O(N__12326),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_7 ));
    InMux I__1040 (
            .O(N__12323),
            .I(N__12320));
    LocalMux I__1039 (
            .O(N__12320),
            .I(N__12317));
    Span4Mux_v I__1038 (
            .O(N__12317),
            .I(N__12314));
    Span4Mux_s1_h I__1037 (
            .O(N__12314),
            .I(N__12311));
    Odrv4 I__1036 (
            .O(N__12311),
            .I(\processor_zipi8.stack_memory_5 ));
    InMux I__1035 (
            .O(N__12308),
            .I(N__12305));
    LocalMux I__1034 (
            .O(N__12305),
            .I(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_5 ));
    CascadeMux I__1033 (
            .O(N__12302),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_5_cascade_ ));
    InMux I__1032 (
            .O(N__12299),
            .I(N__12296));
    LocalMux I__1031 (
            .O(N__12296),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_5 ));
    CascadeMux I__1030 (
            .O(N__12293),
            .I(\processor_zipi8.port_id_5_cascade_ ));
    InMux I__1029 (
            .O(N__12290),
            .I(N__12287));
    LocalMux I__1028 (
            .O(N__12287),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_5 ));
    CascadeMux I__1027 (
            .O(N__12284),
            .I(N__12280));
    CascadeMux I__1026 (
            .O(N__12283),
            .I(N__12277));
    InMux I__1025 (
            .O(N__12280),
            .I(N__12274));
    InMux I__1024 (
            .O(N__12277),
            .I(N__12271));
    LocalMux I__1023 (
            .O(N__12274),
            .I(N__12268));
    LocalMux I__1022 (
            .O(N__12271),
            .I(N__12265));
    Span4Mux_v I__1021 (
            .O(N__12268),
            .I(N__12259));
    Span4Mux_h I__1020 (
            .O(N__12265),
            .I(N__12256));
    InMux I__1019 (
            .O(N__12264),
            .I(N__12249));
    InMux I__1018 (
            .O(N__12263),
            .I(N__12249));
    InMux I__1017 (
            .O(N__12262),
            .I(N__12249));
    Odrv4 I__1016 (
            .O(N__12259),
            .I(\processor_zipi8.port_id_5 ));
    Odrv4 I__1015 (
            .O(N__12256),
            .I(\processor_zipi8.port_id_5 ));
    LocalMux I__1014 (
            .O(N__12249),
            .I(\processor_zipi8.port_id_5 ));
    InMux I__1013 (
            .O(N__12242),
            .I(N__12239));
    LocalMux I__1012 (
            .O(N__12239),
            .I(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_5 ));
    InMux I__1011 (
            .O(N__12236),
            .I(N__12233));
    LocalMux I__1010 (
            .O(N__12233),
            .I(N__12230));
    Odrv4 I__1009 (
            .O(N__12230),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI88F42_7 ));
    CascadeMux I__1008 (
            .O(N__12227),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV3DI8_7_cascade_ ));
    CascadeMux I__1007 (
            .O(N__12224),
            .I(N__12221));
    InMux I__1006 (
            .O(N__12221),
            .I(N__12218));
    LocalMux I__1005 (
            .O(N__12218),
            .I(N__12215));
    Odrv12 I__1004 (
            .O(N__12215),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIM5NP1_7 ));
    InMux I__1003 (
            .O(N__12212),
            .I(N__12209));
    LocalMux I__1002 (
            .O(N__12209),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_7 ));
    InMux I__1001 (
            .O(N__12206),
            .I(N__12203));
    LocalMux I__1000 (
            .O(N__12203),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINR4G8_7 ));
    CascadeMux I__999 (
            .O(N__12200),
            .I(\processor_zipi8.port_id_7_cascade_ ));
    CascadeMux I__998 (
            .O(N__12197),
            .I(N__12193));
    CascadeMux I__997 (
            .O(N__12196),
            .I(N__12190));
    InMux I__996 (
            .O(N__12193),
            .I(N__12187));
    InMux I__995 (
            .O(N__12190),
            .I(N__12184));
    LocalMux I__994 (
            .O(N__12187),
            .I(N__12181));
    LocalMux I__993 (
            .O(N__12184),
            .I(N__12178));
    Span4Mux_v I__992 (
            .O(N__12181),
            .I(N__12172));
    Span4Mux_h I__991 (
            .O(N__12178),
            .I(N__12169));
    InMux I__990 (
            .O(N__12177),
            .I(N__12162));
    InMux I__989 (
            .O(N__12176),
            .I(N__12162));
    InMux I__988 (
            .O(N__12175),
            .I(N__12162));
    Odrv4 I__987 (
            .O(N__12172),
            .I(\processor_zipi8.port_id_7 ));
    Odrv4 I__986 (
            .O(N__12169),
            .I(\processor_zipi8.port_id_7 ));
    LocalMux I__985 (
            .O(N__12162),
            .I(\processor_zipi8.port_id_7 ));
    CascadeMux I__984 (
            .O(N__12155),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_5_cascade_ ));
    CascadeMux I__983 (
            .O(N__12152),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_5_cascade_ ));
    CascadeMux I__982 (
            .O(N__12149),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_5_cascade_ ));
    InMux I__981 (
            .O(N__12146),
            .I(N__12143));
    LocalMux I__980 (
            .O(N__12143),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_5 ));
    CascadeMux I__979 (
            .O(N__12140),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_5_cascade_ ));
    InMux I__978 (
            .O(N__12137),
            .I(N__12134));
    LocalMux I__977 (
            .O(N__12134),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_5 ));
    CascadeMux I__976 (
            .O(N__12131),
            .I(\processor_zipi8.flags_i.un5_shift_carry_value_cascade_ ));
    CascadeMux I__975 (
            .O(N__12128),
            .I(\processor_zipi8.flags_i.shift_carry_value_1_0_0_cascade_ ));
    InMux I__974 (
            .O(N__12125),
            .I(N__12122));
    LocalMux I__973 (
            .O(N__12122),
            .I(N__12119));
    Span4Mux_v I__972 (
            .O(N__12119),
            .I(N__12116));
    Odrv4 I__971 (
            .O(N__12116),
            .I(\processor_zipi8.stack_i.data_out_ram_0 ));
    InMux I__970 (
            .O(N__12113),
            .I(N__12110));
    LocalMux I__969 (
            .O(N__12110),
            .I(\processor_zipi8.shadow_carry_flag ));
    CascadeMux I__968 (
            .O(N__12107),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_7_cascade_ ));
    InMux I__967 (
            .O(N__12104),
            .I(N__12098));
    InMux I__966 (
            .O(N__12103),
            .I(N__12098));
    LocalMux I__965 (
            .O(N__12098),
            .I(N__12095));
    Span4Mux_v I__964 (
            .O(N__12095),
            .I(N__12092));
    Odrv4 I__963 (
            .O(N__12092),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_7 ));
    InMux I__962 (
            .O(N__12089),
            .I(N__12086));
    LocalMux I__961 (
            .O(N__12086),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_7 ));
    CascadeMux I__960 (
            .O(N__12083),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_7_cascade_ ));
    CascadeMux I__959 (
            .O(N__12080),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_7_cascade_ ));
    InMux I__958 (
            .O(N__12077),
            .I(N__12074));
    LocalMux I__957 (
            .O(N__12074),
            .I(N__12071));
    Span4Mux_s1_h I__956 (
            .O(N__12071),
            .I(N__12068));
    Odrv4 I__955 (
            .O(N__12068),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_7 ));
    InMux I__954 (
            .O(N__12065),
            .I(N__12062));
    LocalMux I__953 (
            .O(N__12062),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_7 ));
    CascadeMux I__952 (
            .O(N__12059),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_7_cascade_ ));
    CascadeMux I__951 (
            .O(N__12056),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_7_cascade_ ));
    InMux I__950 (
            .O(N__12053),
            .I(N__12050));
    LocalMux I__949 (
            .O(N__12050),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_7 ));
    CascadeMux I__948 (
            .O(N__12047),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_7_cascade_ ));
    CascadeMux I__947 (
            .O(N__12044),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_7_cascade_ ));
    InMux I__946 (
            .O(N__12041),
            .I(N__12035));
    InMux I__945 (
            .O(N__12040),
            .I(N__12035));
    LocalMux I__944 (
            .O(N__12035),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_7 ));
    CascadeMux I__943 (
            .O(N__12032),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_7_cascade_ ));
    InMux I__942 (
            .O(N__12029),
            .I(N__12023));
    InMux I__941 (
            .O(N__12028),
            .I(N__12023));
    LocalMux I__940 (
            .O(N__12023),
            .I(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_7 ));
    ICE_GB \processor_zipi8.state_machine_i.t_state_RNIA073_2  (
            .USERSIGNALTOGLOBALBUFFER(N__13448),
            .GLOBALBUFFEROUTPUT(bram_enable_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__7_LC_1_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__7_LC_1_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__7_LC_1_2_0 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__7_LC_1_2_0  (
            .in0(N__33312),
            .in1(N__32974),
            .in2(N__36522),
            .in3(N__34765),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33634),
            .ce(N__14864),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_7_LC_1_3_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_7_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_7_LC_1_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_7_LC_1_3_3  (
            .in0(N__37469),
            .in1(N__16426),
            .in2(_gnd_net_),
            .in3(N__13102),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__6_LC_1_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__6_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__6_LC_1_4_0 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__6_LC_1_4_0  (
            .in0(N__34084),
            .in1(N__29265),
            .in2(N__36701),
            .in3(N__29707),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33623),
            .ce(N__25944),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__7_LC_1_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__7_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__7_LC_1_4_1 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__7_LC_1_4_1  (
            .in0(N__32973),
            .in1(N__34085),
            .in2(N__36700),
            .in3(N__33340),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33623),
            .ce(N__25944),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_7_LC_1_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_7_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_7_LC_1_5_0 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_7_LC_1_5_0  (
            .in0(N__34079),
            .in1(N__32824),
            .in2(N__33320),
            .in3(N__36050),
            .lcout(\processor_zipi8.alu_result_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__7_LC_1_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__7_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__7_LC_1_5_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__7_LC_1_5_1  (
            .in0(N__36051),
            .in1(N__33270),
            .in2(N__32898),
            .in3(N__34080),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33614),
            .ce(N__25339),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_7_LC_1_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_7_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_7_LC_1_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_7_LC_1_5_2  (
            .in0(N__12028),
            .in1(N__13150),
            .in2(_gnd_net_),
            .in3(N__37498),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_7_LC_1_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_7_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_7_LC_1_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_7_LC_1_5_3  (
            .in0(N__37499),
            .in1(N__23782),
            .in2(_gnd_net_),
            .in3(N__12040),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_7_LC_1_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_7_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_7_LC_1_5_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_7_LC_1_5_4  (
            .in0(N__12053),
            .in1(N__28653),
            .in2(N__12047),
            .in3(N__29013),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_7_LC_1_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_7_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_7_LC_1_5_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_7_LC_1_5_5  (
            .in0(N__28654),
            .in1(N__20411),
            .in2(N__12044),
            .in3(N__20453),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIP1UE1_7_LC_1_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIP1UE1_7_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIP1UE1_7_LC_1_5_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIP1UE1_7_LC_1_5_6  (
            .in0(N__12041),
            .in1(N__31699),
            .in2(N__23786),
            .in3(N__30993),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI88F42_7_LC_1_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI88F42_7_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI88F42_7_LC_1_5_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI88F42_7_LC_1_5_7  (
            .in0(N__31700),
            .in1(N__13151),
            .in2(N__12032),
            .in3(N__12029),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI88F42_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_7_LC_1_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_7_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_7_LC_1_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_7_LC_1_6_0  (
            .in0(N__13300),
            .in1(N__12103),
            .in2(_gnd_net_),
            .in3(N__37496),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI92021_7_LC_1_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI92021_7_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI92021_7_LC_1_6_1 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI92021_7_LC_1_6_1  (
            .in0(N__13202),
            .in1(N__31702),
            .in2(N__31016),
            .in3(N__16469),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIM5NP1_7_LC_1_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIM5NP1_7_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIM5NP1_7_LC_1_6_2 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIM5NP1_7_LC_1_6_2  (
            .in0(N__13301),
            .in1(N__31750),
            .in2(N__12107),
            .in3(N__12104),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIM5NP1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_7_LC_1_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_7_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_7_LC_1_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_7_LC_1_6_3  (
            .in0(N__37497),
            .in1(N__16468),
            .in2(_gnd_net_),
            .in3(N__13201),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_7_LC_1_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_7_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_7_LC_1_6_4 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_7_LC_1_6_4  (
            .in0(N__29005),
            .in1(N__12089),
            .in2(N__12083),
            .in3(N__28655),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_7_LC_1_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_7_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_7_LC_1_6_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_7_LC_1_6_5  (
            .in0(N__28656),
            .in1(N__13232),
            .in2(N__12080),
            .in3(N__12077),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_7_LC_1_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_7_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_7_LC_1_6_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_7_LC_1_6_6  (
            .in0(N__12065),
            .in1(N__25669),
            .in2(N__12059),
            .in3(N__25792),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_7_LC_1_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_7_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_7_LC_1_6_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_7_LC_1_6_7  (
            .in0(N__25670),
            .in1(N__28310),
            .in2(N__12056),
            .in3(N__20933),
            .lcout(\processor_zipi8.sy_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_5_LC_1_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_5_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_5_LC_1_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_5_LC_1_7_0  (
            .in0(N__13324),
            .in1(N__13279),
            .in2(_gnd_net_),
            .in3(N__37494),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI5UV11_5_LC_1_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI5UV11_5_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI5UV11_5_LC_1_7_1 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI5UV11_5_LC_1_7_1  (
            .in0(N__13223),
            .in1(N__31696),
            .in2(N__31015),
            .in3(N__16496),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIETMP1_5_LC_1_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIETMP1_5_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIETMP1_5_LC_1_7_2 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIETMP1_5_LC_1_7_2  (
            .in0(N__13325),
            .in1(N__31697),
            .in2(N__12155),
            .in3(N__13280),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_5_LC_1_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_5_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_5_LC_1_7_3 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_5_LC_1_7_3  (
            .in0(N__18104),
            .in1(N__12137),
            .in2(N__13271),
            .in3(N__28622),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_5_LC_1_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_5_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_5_LC_1_7_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_5_LC_1_7_4  (
            .in0(N__24986),
            .in1(N__25660),
            .in2(N__12152),
            .in3(N__25761),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_5_LC_1_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_5_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_5_LC_1_7_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_5_LC_1_7_5  (
            .in0(N__25661),
            .in1(N__22697),
            .in2(N__12149),
            .in3(N__20399),
            .lcout(\processor_zipi8.sy_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_5_LC_1_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_5_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_5_LC_1_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_5_LC_1_7_6  (
            .in0(N__16495),
            .in1(N__13222),
            .in2(_gnd_net_),
            .in3(N__37495),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_5_LC_1_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_5_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_5_LC_1_7_7 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_5_LC_1_7_7  (
            .in0(N__12146),
            .in1(N__28621),
            .in2(N__12140),
            .in3(N__29004),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.shift_carry_RNO_1_LC_1_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.shift_carry_RNO_1_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.shift_carry_RNO_1_LC_1_8_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \processor_zipi8.flags_i.shift_carry_RNO_1_LC_1_8_0  (
            .in0(N__16679),
            .in1(N__17102),
            .in2(_gnd_net_),
            .in3(N__24316),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.un5_shift_carry_value_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.shift_carry_RNO_0_LC_1_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.shift_carry_RNO_0_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.shift_carry_RNO_0_LC_1_8_1 .LUT_INIT=16'b0000010000000111;
    LogicCell40 \processor_zipi8.flags_i.shift_carry_RNO_0_LC_1_8_1  (
            .in0(N__25783),
            .in1(N__24318),
            .in2(N__12131),
            .in3(N__12113),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.shift_carry_value_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.shift_carry_LC_1_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.shift_carry_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.flags_i.shift_carry_LC_1_8_2 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \processor_zipi8.flags_i.shift_carry_LC_1_8_2  (
            .in0(N__17121),
            .in1(N__24317),
            .in2(N__12128),
            .in3(N__21113),
            .lcout(\processor_zipi8.flags_i.shift_carryZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33606),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.shadow_carry_flag_0_LC_1_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_0_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_0_LC_1_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.stack_i.shadow_carry_flag_0_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12125),
            .lcout(\processor_zipi8.shadow_carry_flag ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33606),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU7BG4_7_LC_1_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU7BG4_7_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU7BG4_7_LC_1_8_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU7BG4_7_LC_1_8_4  (
            .in0(N__12236),
            .in1(N__27439),
            .in2(N__20252),
            .in3(N__27636),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV3DI8_7_LC_1_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV3DI8_7_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV3DI8_7_LC_1_8_5 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV3DI8_7_LC_1_8_5  (
            .in0(N__27441),
            .in1(N__28259),
            .in2(N__22883),
            .in3(N__20222),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV3DI8_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5S0IH_7_LC_1_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5S0IH_7_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5S0IH_7_LC_1_8_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5S0IH_7_LC_1_8_6  (
            .in0(N__12206),
            .in1(_gnd_net_),
            .in2(N__12227),
            .in3(N__22233),
            .lcout(\processor_zipi8.sx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINR4G8_7_LC_1_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINR4G8_7_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINR4G8_7_LC_1_8_7 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINR4G8_7_LC_1_8_7  (
            .in0(N__27440),
            .in1(N__13115),
            .in2(N__12224),
            .in3(N__12212),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINR4G8_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_7_LC_1_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_7_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_7_LC_1_9_0 .LUT_INIT=16'b0101011111110111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_7_LC_1_9_0  (
            .in0(N__12176),
            .in1(N__19588),
            .in2(N__16684),
            .in3(N__19639),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_0_LC_1_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_0_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_0_LC_1_9_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_0_LC_1_9_1  (
            .in0(N__12368),
            .in1(N__21447),
            .in2(_gnd_net_),
            .in3(N__25782),
            .lcout(\processor_zipi8.port_id_7 ),
            .ltout(\processor_zipi8.port_id_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_7_LC_1_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_7_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_7_LC_1_9_2 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_7_LC_1_9_2  (
            .in0(N__16667),
            .in1(N__19208),
            .in2(N__12200),
            .in3(N__19589),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_7_LC_1_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_7_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_7_LC_1_9_3 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_7_LC_1_9_3  (
            .in0(N__19207),
            .in1(N__12177),
            .in2(N__16683),
            .in3(N__24013),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_7_LC_1_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_7_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_7_LC_1_9_4 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_7_LC_1_9_4  (
            .in0(N__12175),
            .in1(N__19486),
            .in2(N__16685),
            .in3(N__19799),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_7_LC_1_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_7_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_7_LC_1_9_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_7_LC_1_9_5  (
            .in0(N__12347),
            .in1(N__12338),
            .in2(N__12332),
            .in3(N__12329),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_5_LC_1_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_5_LC_1_9_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_5_LC_1_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_5_LC_1_9_6  (
            .in0(N__12323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33608),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNID2G21_5_LC_1_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNID2G21_5_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNID2G21_5_LC_1_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNID2G21_5_LC_1_9_7  (
            .in0(N__29015),
            .in1(N__12308),
            .in2(_gnd_net_),
            .in3(N__21446),
            .lcout(\processor_zipi8.pc_vector_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_5_LC_1_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_5_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_5_LC_1_10_0 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_5_LC_1_10_0  (
            .in0(N__12262),
            .in1(N__19478),
            .in2(N__18784),
            .in3(N__19797),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_5_LC_1_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_5_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_5_LC_1_10_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_5_LC_1_10_1  (
            .in0(N__12242),
            .in1(N__12290),
            .in2(N__12302),
            .in3(N__12299),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_5_LC_1_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_5_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_5_LC_1_10_2 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_5_LC_1_10_2  (
            .in0(N__12263),
            .in1(N__19580),
            .in2(N__18783),
            .in3(N__19201),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_2_0_LC_1_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_2_0_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_2_0_LC_1_10_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_2_0_LC_1_10_3  (
            .in0(N__12383),
            .in1(N__21452),
            .in2(_gnd_net_),
            .in3(N__29014),
            .lcout(\processor_zipi8.port_id_5 ),
            .ltout(\processor_zipi8.port_id_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_5_LC_1_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_5_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_5_LC_1_10_4 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_5_LC_1_10_4  (
            .in0(N__18765),
            .in1(N__19579),
            .in2(N__12293),
            .in3(N__19632),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_5_LC_1_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_5_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_5_LC_1_10_5 .LUT_INIT=16'b1111111101000111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_5_LC_1_10_5  (
            .in0(N__19200),
            .in1(N__12264),
            .in2(N__24014),
            .in3(N__18766),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_9_LC_1_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_9_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_9_LC_1_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_9_LC_1_10_6  (
            .in0(N__12437),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33609),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_4_LC_1_10_7 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_4_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_4_LC_1_10_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_4_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__12428),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33609),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIG4G21_7_LC_1_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIG4G21_7_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIG4G21_7_LC_1_11_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIG4G21_7_LC_1_11_0  (
            .in0(N__13865),
            .in1(N__21453),
            .in2(_gnd_net_),
            .in3(N__25784),
            .lcout(\processor_zipi8.pc_vector_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_8_LC_1_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_8_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_8_LC_1_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_8_LC_1_11_1  (
            .in0(N__12419),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33613),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_10_LC_1_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_10_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_10_LC_1_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_10_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12407),
            .lcout(\processor_zipi8.return_vector_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33613),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIJ6G21_9_LC_1_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIJ6G21_9_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIJ6G21_9_LC_1_12_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIJ6G21_9_LC_1_12_0  (
            .in0(N__12395),
            .in1(N__21455),
            .in2(_gnd_net_),
            .in3(N__31694),
            .lcout(\processor_zipi8.pc_vector_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNING29O_5_LC_1_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNING29O_5_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNING29O_5_LC_1_12_1 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNING29O_5_LC_1_12_1  (
            .in0(N__12382),
            .in1(N__17882),
            .in2(N__13940),
            .in3(N__17800),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIOI39O_6_LC_1_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIOI39O_6_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIOI39O_6_LC_1_12_2 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIOI39O_6_LC_1_12_2  (
            .in0(N__17801),
            .in1(N__13730),
            .in2(N__17890),
            .in3(N__13406),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIPK49O_7_LC_1_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIPK49O_7_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIPK49O_7_LC_1_12_3 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIPK49O_7_LC_1_12_3  (
            .in0(N__12367),
            .in1(N__17886),
            .in2(N__14123),
            .in3(N__17802),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNII5G21_8_LC_1_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNII5G21_8_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNII5G21_8_LC_1_12_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNII5G21_8_LC_1_12_4  (
            .in0(N__12803),
            .in1(N__21454),
            .in2(_gnd_net_),
            .in3(N__31021),
            .lcout(\processor_zipi8.pc_vector_8 ),
            .ltout(\processor_zipi8.pc_vector_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_8_LC_1_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_8_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_8_LC_1_12_5 .LUT_INIT=16'b0011100110011001;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_8_LC_1_12_5  (
            .in0(N__12878),
            .in1(N__12443),
            .in2(N__12797),
            .in3(N__15939),
            .lcout(address_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33622),
            .ce(N__15763),
            .sr(N__17401));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI9LLGO_9_LC_1_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI9LLGO_9_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI9LLGO_9_LC_1_12_6 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNI9LLGO_9_LC_1_12_6  (
            .in0(N__17803),
            .in1(N__12678),
            .in2(N__17891),
            .in3(N__21706),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_9 ),
            .ltout(\processor_zipi8.program_counter_i.half_pc_0_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_9_LC_1_12_7 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_9_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_9_LC_1_12_7 .LUT_INIT=16'b0111000010001111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_9_LC_1_12_7  (
            .in0(N__14380),
            .in1(N__15940),
            .in2(N__12794),
            .in3(N__14366),
            .lcout(address_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33622),
            .ce(N__15763),
            .sr(N__17401));
    defparam \processor_zipi8.program_counter_i.pc_RNIDL1F5_10_LC_1_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_RNIDL1F5_10_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_RNIDL1F5_10_LC_1_13_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_RNIDL1F5_10_LC_1_13_0  (
            .in0(N__17776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12498),
            .lcout(),
            .ltout(\processor_zipi8.program_counter_i.un380_half_pc_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_RNIDJA501_10_LC_1_13_1 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_RNIDJA501_10_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_RNIDJA501_10_LC_1_13_1 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_RNIDJA501_10_LC_1_13_1  (
            .in0(N__17861),
            .in1(N__22013),
            .in2(N__12635),
            .in3(N__12449),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_10 ),
            .ltout(\processor_zipi8.program_counter_i.half_pc_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_10_LC_1_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_10_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_10_LC_1_13_2 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \processor_zipi8.program_counter_i.pc_10_LC_1_13_2  (
            .in0(N__19058),
            .in1(N__12499),
            .in2(N__12632),
            .in3(N__14354),
            .lcout(address_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33626),
            .ce(),
            .sr(N__17429));
    defparam \processor_zipi8.program_counter_i.un395_half_pc_LC_1_13_3 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.un395_half_pc_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.un395_half_pc_LC_1_13_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \processor_zipi8.program_counter_i.un395_half_pc_LC_1_13_3  (
            .in0(N__15937),
            .in1(N__21456),
            .in2(N__12464),
            .in3(N__27641),
            .lcout(\processor_zipi8.program_counter_i.un395_half_pcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIQQO068_7_LC_1_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIQQO068_7_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIQQO068_7_LC_1_13_4 .LUT_INIT=16'b1101010100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIQQO068_7_LC_1_13_4  (
            .in0(N__14236),
            .in1(N__15935),
            .in2(N__14261),
            .in3(N__14267),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_46_7 ),
            .ltout(\processor_zipi8.program_counter_i.carry_pc_46_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIT0QD69_8_LC_1_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIT0QD69_8_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIT0QD69_8_LC_1_13_5 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIT0QD69_8_LC_1_13_5  (
            .in0(N__15936),
            .in1(N__13049),
            .in2(N__13040),
            .in3(N__12874),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_52_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8JKGO_8_LC_1_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8JKGO_8_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8JKGO_8_LC_1_13_6 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNI8JKGO_8_LC_1_13_6  (
            .in0(N__17775),
            .in1(N__17860),
            .in2(N__12943),
            .in3(N__21111),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNO_0_LC_1_14_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_0_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_0_LC_1_14_0 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNO_0_LC_1_14_0  (
            .in0(N__16889),
            .in1(N__12836),
            .in2(N__12860),
            .in3(N__17903),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.zero_flag_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_LC_1_14_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_LC_1_14_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.flags_i.zero_flag_LC_1_14_1 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_LC_1_14_1  (
            .in0(N__17400),
            .in1(N__17506),
            .in2(N__12863),
            .in3(N__18033),
            .lcout(\processor_zipi8.zero_flag ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33633),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.shadow_zero_flag_LC_1_14_2 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.shadow_zero_flag_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.shadow_zero_flag_LC_1_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.stack_i.shadow_zero_flag_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12809),
            .lcout(\processor_zipi8.shadow_zero_flag ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33633),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_6_LC_1_14_3 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_6_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_6_LC_1_14_3 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_6_LC_1_14_3  (
            .in0(N__34083),
            .in1(N__29371),
            .in2(N__29736),
            .in3(N__35861),
            .lcout(),
            .ltout(\processor_zipi8.alu_result_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNO_1_LC_1_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_1_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_1_LC_1_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNO_1_LC_1_14_4  (
            .in0(N__12851),
            .in1(N__12830),
            .in2(N__12839),
            .in3(N__13091),
            .lcout(\processor_zipi8.flags_i.zero_flag_3_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_5_LC_1_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_5_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_5_LC_1_14_5 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_5_LC_1_14_5  (
            .in0(N__34081),
            .in1(N__29952),
            .in2(N__30492),
            .in3(N__35859),
            .lcout(\processor_zipi8.alu_result_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.shadow_carry_flag_1_LC_1_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_1_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_1_LC_1_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.stack_i.shadow_carry_flag_1_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12824),
            .lcout(\processor_zipi8.stack_i.shadow_zero_value ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33633),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_3_LC_1_14_7 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_3_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_3_LC_1_14_7 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_3_LC_1_14_7  (
            .in0(N__34082),
            .in1(N__37628),
            .in2(N__38174),
            .in3(N__35860),
            .lcout(\processor_zipi8.alu_result_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI0LOT3_LC_1_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI0LOT3_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI0LOT3_LC_1_15_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI0LOT3_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__14658),
            .in2(_gnd_net_),
            .in3(N__14325),
            .lcout(\processor_zipi8.flags_i.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNICAJR_LC_1_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNICAJR_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNICAJR_LC_1_15_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNICAJR_LC_1_15_1  (
            .in0(N__18029),
            .in1(N__17989),
            .in2(_gnd_net_),
            .in3(N__24112),
            .lcout(\processor_zipi8.flags_i.m49_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIJK644_LC_1_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIJK644_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIJK644_LC_1_15_3 .LUT_INIT=16'b0011011100001000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIJK644_LC_1_15_3  (
            .in0(N__14327),
            .in1(N__19042),
            .in2(N__16290),
            .in3(N__14660),
            .lcout(\processor_zipi8.flags_i.m82_1 ),
            .ltout(\processor_zipi8.flags_i.m82_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.stack_pointer_1_LC_1_15_4 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.stack_pointer_1_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.stack_pointer_1_LC_1_15_4 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \processor_zipi8.stack_i.stack_pointer_1_LC_1_15_4  (
            .in0(N__14560),
            .in1(N__17394),
            .in2(N__13085),
            .in3(N__16276),
            .lcout(\processor_zipi8.stack_pointer_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33641),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIJSPM4_LC_1_15_5 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIJSPM4_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIJSPM4_LC_1_15_5 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIJSPM4_LC_1_15_5  (
            .in0(N__16275),
            .in1(N__13082),
            .in2(N__17416),
            .in3(N__14559),
            .lcout(\processor_zipi8.zero_flag_RNIJSPM4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIALV04_LC_1_15_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIALV04_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIALV04_LC_1_15_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIALV04_LC_1_15_6  (
            .in0(N__14659),
            .in1(N__16271),
            .in2(_gnd_net_),
            .in3(N__14326),
            .lcout(\processor_zipi8.flags_i.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI6N578_LC_1_16_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI6N578_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI6N578_LC_1_16_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI6N578_LC_1_16_3  (
            .in0(N__14486),
            .in1(N__14455),
            .in2(N__15167),
            .in3(N__13058),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.m61_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNID5QI8_LC_1_16_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNID5QI8_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNID5QI8_LC_1_16_4 .LUT_INIT=16'b0010001101100101;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNID5QI8_LC_1_16_4  (
            .in0(N__15165),
            .in1(N__17260),
            .in2(N__13052),
            .in3(N__16280),
            .lcout(\processor_zipi8.flags_i.i14_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI3VC94_LC_1_16_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI3VC94_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI3VC94_LC_1_16_6 .LUT_INIT=16'b0011101000110101;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI3VC94_LC_1_16_6  (
            .in0(N__14456),
            .in1(N__14661),
            .in2(N__16291),
            .in3(N__14487),
            .lcout(\processor_zipi8.flags_i.zero_flag_RNI3VCZ0Z94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__7_LC_2_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__7_LC_2_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__7_LC_2_2_0 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__7_LC_2_2_0  (
            .in0(N__34520),
            .in1(N__36661),
            .in2(N__33013),
            .in3(N__33316),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33642),
            .ce(N__26167),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNITSK21_6_LC_2_3_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNITSK21_6_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNITSK21_6_LC_2_3_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNITSK21_6_LC_2_3_0  (
            .in0(N__13130),
            .in1(N__31745),
            .in2(N__16445),
            .in3(N__30985),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIGUSR1_6_LC_2_3_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIGUSR1_6_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIGUSR1_6_LC_2_3_1 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIGUSR1_6_LC_2_3_1  (
            .in0(N__13262),
            .in1(N__31744),
            .in2(N__13133),
            .in3(N__16394),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIGUSR1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_6_LC_2_3_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_6_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_6_LC_2_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_6_LC_2_3_2  (
            .in0(N__16441),
            .in1(N__13129),
            .in2(_gnd_net_),
            .in3(N__37468),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__6_LC_2_3_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__6_LC_2_3_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__6_LC_2_3_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__6_LC_2_3_3  (
            .in0(N__34303),
            .in1(N__36557),
            .in2(N__29365),
            .in3(N__29706),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33636),
            .ce(N__18076),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_6_LC_2_3_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_6_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_6_LC_2_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_6_LC_2_3_4  (
            .in0(N__16393),
            .in1(N__13261),
            .in2(_gnd_net_),
            .in3(N__37467),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIVUK21_7_LC_2_3_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIVUK21_7_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIVUK21_7_LC_2_3_5 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIVUK21_7_LC_2_3_5  (
            .in0(N__30986),
            .in1(N__16427),
            .in2(N__31751),
            .in3(N__13103),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIK2TR1_7_LC_2_3_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIK2TR1_7_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIK2TR1_7_LC_2_3_6 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIK2TR1_7_LC_2_3_6  (
            .in0(N__13250),
            .in1(N__16541),
            .in2(N__13118),
            .in3(N__31749),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIK2TR1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__7_LC_2_3_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__7_LC_2_3_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__7_LC_2_3_7 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__7_LC_2_3_7  (
            .in0(N__34304),
            .in1(N__32978),
            .in2(N__33359),
            .in3(N__36558),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33636),
            .ce(N__18076),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_6_LC_2_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_6_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_6_LC_2_4_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_6_LC_2_4_0  (
            .in0(N__13210),
            .in1(N__37394),
            .in2(_gnd_net_),
            .in3(N__16483),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI70021_6_LC_2_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI70021_6_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI70021_6_LC_2_4_1 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI70021_6_LC_2_4_1  (
            .in0(N__16484),
            .in1(N__31698),
            .in2(N__31014),
            .in3(N__13211),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNII1NP1_6_LC_2_4_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNII1NP1_6_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNII1NP1_6_LC_2_4_2 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNII1NP1_6_LC_2_4_2  (
            .in0(N__13430),
            .in1(N__31701),
            .in2(N__13190),
            .in3(N__13316),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNII1NP1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_6_LC_2_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_6_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_6_LC_2_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_6_LC_2_4_3  (
            .in0(N__37395),
            .in1(N__13315),
            .in2(_gnd_net_),
            .in3(N__13429),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_6_LC_2_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_6_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_6_LC_2_4_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_6_LC_2_4_4  (
            .in0(N__13187),
            .in1(N__28649),
            .in2(N__13181),
            .in3(N__29012),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_6_LC_2_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_6_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_6_LC_2_4_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_6_LC_2_4_5  (
            .in0(N__28650),
            .in1(N__13178),
            .in2(N__13169),
            .in3(N__13166),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_6_LC_2_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_6_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_6_LC_2_4_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_6_LC_2_4_6  (
            .in0(N__14753),
            .in1(N__25667),
            .in2(N__13157),
            .in3(N__25785),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_6_LC_2_4_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_6_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_6_LC_2_4_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_6_LC_2_4_7  (
            .in0(N__25668),
            .in1(N__23828),
            .in2(N__13154),
            .in3(N__24611),
            .lcout(\processor_zipi8.sy_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__0_LC_2_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__0_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__0_LC_2_5_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__0_LC_2_5_0  (
            .in0(N__34751),
            .in1(N__36553),
            .in2(N__32460),
            .in3(N__32026),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__1_LC_2_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__1_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__1_LC_2_5_1 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__1_LC_2_5_1  (
            .in0(N__36549),
            .in1(N__34756),
            .in2(N__39233),
            .in3(N__39592),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__2_LC_2_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__2_LC_2_5_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__2_LC_2_5_2 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__2_LC_2_5_2  (
            .in0(N__38556),
            .in1(N__36554),
            .in2(N__34840),
            .in3(N__38730),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__3_LC_2_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__3_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__3_LC_2_5_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__3_LC_2_5_3  (
            .in0(N__36550),
            .in1(N__34754),
            .in2(N__38184),
            .in3(N__37825),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__4_LC_2_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__4_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__4_LC_2_5_4 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__4_LC_2_5_4  (
            .in0(N__34752),
            .in1(N__36555),
            .in2(N__35560),
            .in3(N__35156),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__5_LC_2_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__5_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__5_LC_2_5_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__5_LC_2_5_5  (
            .in0(N__36551),
            .in1(N__34755),
            .in2(N__30499),
            .in3(N__29951),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__6_LC_2_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__6_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__6_LC_2_5_6 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__6_LC_2_5_6  (
            .in0(N__34753),
            .in1(N__36556),
            .in2(N__29705),
            .in3(N__29315),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__7_LC_2_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__7_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__7_LC_2_5_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram8__7_LC_2_5_7  (
            .in0(N__36552),
            .in1(N__33271),
            .in2(N__32995),
            .in3(N__34760),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram8_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33625),
            .ce(N__14876),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__0_LC_2_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__0_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__0_LC_2_6_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__0_LC_2_6_0  (
            .in0(N__34556),
            .in1(N__36596),
            .in2(N__32433),
            .in3(N__32025),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33616),
            .ce(N__20288),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__2_LC_2_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__2_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__2_LC_2_6_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__2_LC_2_6_1  (
            .in0(N__36593),
            .in1(N__34558),
            .in2(N__38802),
            .in3(N__38557),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33616),
            .ce(N__20288),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__3_LC_2_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__3_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__3_LC_2_6_2 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__3_LC_2_6_2  (
            .in0(N__37774),
            .in1(N__38154),
            .in2(N__34764),
            .in3(N__36598),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33616),
            .ce(N__20288),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__5_LC_2_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__5_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__5_LC_2_6_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__5_LC_2_6_3  (
            .in0(N__36594),
            .in1(N__34559),
            .in2(N__30508),
            .in3(N__29950),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33616),
            .ce(N__20288),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_5_LC_2_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_5_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_5_LC_2_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_5_LC_2_6_4  (
            .in0(N__18296),
            .in1(N__18274),
            .in2(_gnd_net_),
            .in3(N__37484),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__6_LC_2_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__6_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__6_LC_2_6_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__6_LC_2_6_5  (
            .in0(N__36595),
            .in1(N__34560),
            .in2(N__29770),
            .in3(N__29316),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33616),
            .ce(N__20288),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__7_LC_2_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__7_LC_2_6_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__7_LC_2_6_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__7_LC_2_6_6  (
            .in0(N__34557),
            .in1(N__36597),
            .in2(N__33017),
            .in3(N__33319),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33616),
            .ce(N__20288),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_7_LC_2_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_7_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_7_LC_2_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_7_LC_2_6_7  (
            .in0(N__37485),
            .in1(N__16537),
            .in2(_gnd_net_),
            .in3(N__13243),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__0_LC_2_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__0_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__0_LC_2_7_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__0_LC_2_7_0  (
            .in0(N__34742),
            .in1(N__36370),
            .in2(N__32432),
            .in3(N__32024),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__1_LC_2_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__1_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__1_LC_2_7_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__1_LC_2_7_1  (
            .in0(N__36366),
            .in1(N__34745),
            .in2(N__39598),
            .in3(N__39224),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__2_LC_2_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__2_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__2_LC_2_7_2 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__2_LC_2_7_2  (
            .in0(N__38513),
            .in1(N__36371),
            .in2(N__34839),
            .in3(N__38729),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__3_LC_2_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__3_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__3_LC_2_7_3 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__3_LC_2_7_3  (
            .in0(N__36367),
            .in1(N__34747),
            .in2(N__37862),
            .in3(N__38147),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__4_LC_2_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__4_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__4_LC_2_7_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__4_LC_2_7_4  (
            .in0(N__34743),
            .in1(N__36372),
            .in2(N__35211),
            .in3(N__35573),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__5_LC_2_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__5_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__5_LC_2_7_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__5_LC_2_7_5  (
            .in0(N__36368),
            .in1(N__34746),
            .in2(N__30444),
            .in3(N__29894),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__6_LC_2_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__6_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__6_LC_2_7_6 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__6_LC_2_7_6  (
            .in0(N__34744),
            .in1(N__29311),
            .in2(N__29769),
            .in3(N__36373),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__7_LC_2_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__7_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__7_LC_2_7_7 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__7_LC_2_7_7  (
            .in0(N__36369),
            .in1(N__33318),
            .in2(N__34841),
            .in3(N__32993),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram11_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33610),
            .ce(N__14897),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__0_LC_2_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__0_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__0_LC_2_8_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__0_LC_2_8_0  (
            .in0(N__34402),
            .in1(N__36201),
            .in2(N__32431),
            .in3(N__32023),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33607),
            .ce(N__14863),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__1_LC_2_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__1_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__1_LC_2_8_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__1_LC_2_8_1  (
            .in0(N__36197),
            .in1(N__39545),
            .in2(N__39228),
            .in3(N__34406),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33607),
            .ce(N__14863),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__2_LC_2_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__2_LC_2_8_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__2_LC_2_8_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__2_LC_2_8_2  (
            .in0(N__34403),
            .in1(N__36202),
            .in2(N__38558),
            .in3(N__38725),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33607),
            .ce(N__14863),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__3_LC_2_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__3_LC_2_8_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__3_LC_2_8_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__3_LC_2_8_3  (
            .in0(N__36198),
            .in1(N__34405),
            .in2(N__38185),
            .in3(N__37797),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33607),
            .ce(N__14863),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_5_LC_2_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_5_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_5_LC_2_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_5_LC_2_8_4  (
            .in0(N__14912),
            .in1(N__13289),
            .in2(_gnd_net_),
            .in3(N__36196),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202 ),
            .ltout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1202_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__5_LC_2_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__5_LC_2_8_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__5_LC_2_8_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__5_LC_2_8_5  (
            .in0(N__36199),
            .in1(N__30461),
            .in2(N__13283),
            .in3(N__34407),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33607),
            .ce(N__14863),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__4_LC_2_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__4_LC_2_8_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__4_LC_2_8_6 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__4_LC_2_8_6  (
            .in0(N__34404),
            .in1(N__35155),
            .in2(N__35569),
            .in3(N__36203),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33607),
            .ce(N__14863),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__6_LC_2_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__6_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__6_LC_2_8_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram10__6_LC_2_8_7  (
            .in0(N__36200),
            .in1(N__29684),
            .in2(N__29366),
            .in3(N__34408),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33607),
            .ce(N__14863),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_6_LC_2_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_6_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_6_LC_2_9_0 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_6_LC_2_9_0  (
            .in0(N__13351),
            .in1(N__19474),
            .in2(N__16633),
            .in3(N__19798),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_6_LC_2_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_6_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_6_LC_2_9_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_6_LC_2_9_1  (
            .in0(N__13331),
            .in1(N__13376),
            .in2(N__13415),
            .in3(N__13412),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_6_LC_2_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_6_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_6_LC_2_9_2 .LUT_INIT=16'b0100111101111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_6_LC_2_9_2  (
            .in0(N__19640),
            .in1(N__16630),
            .in2(N__13362),
            .in3(N__19587),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_1_0_LC_2_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_1_0_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_1_0_LC_2_9_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_1_0_LC_2_9_3  (
            .in0(N__28652),
            .in1(_gnd_net_),
            .in2(N__21458),
            .in3(N__13405),
            .lcout(\processor_zipi8.port_id_6 ),
            .ltout(\processor_zipi8.port_id_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_6_LC_2_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_6_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_6_LC_2_9_4 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_6_LC_2_9_4  (
            .in0(N__16623),
            .in1(N__19586),
            .in2(N__13379),
            .in3(N__19206),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_6_LC_2_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_6_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_6_LC_2_9_5 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_6_LC_2_9_5  (
            .in0(N__19205),
            .in1(N__13355),
            .in2(N__16634),
            .in3(N__24012),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIF3G21_6_LC_2_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIF3G21_6_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIF3G21_6_LC_2_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIF3G21_6_LC_2_9_6  (
            .in0(N__13520),
            .in1(N__21448),
            .in2(_gnd_net_),
            .in3(N__28651),
            .lcout(\processor_zipi8.pc_vector_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_6_LC_2_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_6_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_6_LC_2_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_6_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13529),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33611),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.state_machine_i.t_state_1_LC_2_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.state_machine_i.t_state_1_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.state_machine_i.t_state_1_LC_2_10_0 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \processor_zipi8.state_machine_i.t_state_1_LC_2_10_0  (
            .in0(N__17339),
            .in1(N__19005),
            .in2(N__13460),
            .in3(N__16289),
            .lcout(\processor_zipi8.t_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33615),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_2_LC_2_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_2_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_2_LC_2_10_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_2_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__16868),
            .in2(_gnd_net_),
            .in3(N__17021),
            .lcout(\processor_zipi8.arith_logical_result_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33615),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m38_LC_2_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m38_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m38_LC_2_10_2 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \processor_zipi8.flags_i.m38_LC_2_10_2  (
            .in0(N__13486),
            .in1(N__13879),
            .in2(_gnd_net_),
            .in3(N__15144),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.N_125_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.state_machine_i.run_LC_2_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.state_machine_i.run_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.state_machine_i.run_LC_2_10_3 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \processor_zipi8.state_machine_i.run_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__13501),
            .in2(N__13511),
            .in3(N__17340),
            .lcout(\processor_zipi8.run ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33615),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.shadow_carry_flag_3_LC_2_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_3_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_3_LC_2_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.stack_i.shadow_carry_flag_3_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13508),
            .lcout(\processor_zipi8.special_bit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33615),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.state_machine_i.internal_reset_LC_2_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.state_machine_i.internal_reset_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.state_machine_i.internal_reset_LC_2_10_5 .LUT_INIT=16'b1111111101110011;
    LogicCell40 \processor_zipi8.state_machine_i.internal_reset_LC_2_10_5  (
            .in0(N__13880),
            .in1(N__13500),
            .in2(N__15158),
            .in3(N__13487),
            .lcout(\processor_zipi8.internal_reset ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33615),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_2_LC_2_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_2_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_2_LC_2_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_2_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13466),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33615),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.state_machine_i.t_state_2_LC_2_10_7 .C_ON=1'b0;
    defparam \processor_zipi8.state_machine_i.t_state_2_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.state_machine_i.t_state_2_LC_2_10_7 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \processor_zipi8.state_machine_i.t_state_2_LC_2_10_7  (
            .in0(N__16288),
            .in1(N__13459),
            .in2(N__19041),
            .in3(N__17341),
            .lcout(\processor_zipi8.state_machine_i.bram_enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33615),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_11_LC_2_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_11_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_11_LC_2_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_11_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13436),
            .lcout(\processor_zipi8.return_vector_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33624),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m36_LC_2_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m36_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m36_LC_2_11_1 .LUT_INIT=16'b0001001111011111;
    LogicCell40 \processor_zipi8.flags_i.m36_LC_2_11_1  (
            .in0(N__17255),
            .in1(N__19000),
            .in2(N__15113),
            .in3(N__16287),
            .lcout(\processor_zipi8.flags_i.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.stack_pointer_4_LC_2_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.stack_pointer_4_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.stack_pointer_4_LC_2_11_2 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \processor_zipi8.stack_i.stack_pointer_4_LC_2_11_2  (
            .in0(N__19001),
            .in1(N__15827),
            .in2(N__17379),
            .in3(N__15803),
            .lcout(\processor_zipi8.stack_pointer_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33624),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_7_LC_2_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_7_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_7_LC_2_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_7_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13871),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33624),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_1_LC_2_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_1_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_1_LC_2_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_1_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13859),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33624),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINQ3G8_5_LC_2_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINQ3G8_5_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINQ3G8_5_LC_2_11_6 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINQ3G8_5_LC_2_11_6  (
            .in0(N__13847),
            .in1(N__23663),
            .in2(N__18263),
            .in3(N__27316),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_195_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5QUHH_5_LC_2_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5QUHH_5_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5QUHH_5_LC_2_11_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5QUHH_5_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__22790),
            .in2(N__13835),
            .in3(N__22232),
            .lcout(\processor_zipi8.sx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_4_LC_2_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_4_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_4_LC_2_12_0 .LUT_INIT=16'b0101100110011001;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_4_LC_2_12_0  (
            .in0(N__15332),
            .in1(N__13535),
            .in2(N__15954),
            .in3(N__21245),
            .lcout(address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33627),
            .ce(N__15762),
            .sr(N__17444));
    defparam \processor_zipi8.program_counter_i.pc_esr_6_LC_2_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_6_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_6_LC_2_12_1 .LUT_INIT=16'b0110101001010101;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_6_LC_2_12_1  (
            .in0(N__14303),
            .in1(N__15933),
            .in2(N__14297),
            .in3(N__14276),
            .lcout(address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33627),
            .ce(N__15762),
            .sr(N__17444));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIJE19O_4_LC_2_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIJE19O_4_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIJE19O_4_LC_2_12_2 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIJE19O_4_LC_2_12_2  (
            .in0(N__17881),
            .in1(N__16948),
            .in2(N__13586),
            .in3(N__17799),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_4 ),
            .ltout(\processor_zipi8.program_counter_i.half_pc_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIBG8G55_4_LC_2_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIBG8G55_4_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIBG8G55_4_LC_2_12_3 .LUT_INIT=16'b1000111100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIBG8G55_4_LC_2_12_3  (
            .in0(N__21244),
            .in1(N__15926),
            .in2(N__14309),
            .in3(N__15331),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_28_4 ),
            .ltout(\processor_zipi8.program_counter_i.carry_pc_28_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIOGNL56_5_LC_2_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIOGNL56_5_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIOGNL56_5_LC_2_12_4 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIOGNL56_5_LC_2_12_4  (
            .in0(N__15927),
            .in1(N__14059),
            .in2(N__14306),
            .in3(N__14074),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_34_5 ),
            .ltout(\processor_zipi8.program_counter_i.carry_pc_34_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8K7R57_6_LC_2_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8K7R57_6_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8K7R57_6_LC_2_12_5 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNI8K7R57_6_LC_2_12_5  (
            .in0(N__14293),
            .in1(N__15928),
            .in2(N__14279),
            .in3(N__14275),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_40_6 ),
            .ltout(\processor_zipi8.program_counter_i.carry_pc_40_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_7_LC_2_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_7_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_7_LC_2_12_6 .LUT_INIT=16'b0111100000001111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_7_LC_2_12_6  (
            .in0(N__15934),
            .in1(N__14260),
            .in2(N__14240),
            .in3(N__14237),
            .lcout(address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33627),
            .ce(N__15762),
            .sr(N__17444));
    defparam \processor_zipi8.program_counter_i.pc_esr_5_LC_2_12_7 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_5_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_5_LC_2_12_7 .LUT_INIT=16'b0010101011010101;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_5_LC_2_12_7  (
            .in0(N__14075),
            .in1(N__15932),
            .in2(N__14063),
            .in3(N__14048),
            .lcout(address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33627),
            .ce(N__15762),
            .sr(N__17444));
    defparam \processor_zipi8.program_counter_i.un3_half_pc_LC_2_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.un3_half_pc_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.un3_half_pc_LC_2_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \processor_zipi8.program_counter_i.un3_half_pc_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__17857),
            .in2(_gnd_net_),
            .in3(N__17771),
            .lcout(\processor_zipi8.program_counter_i.un3_half_pcZ0 ),
            .ltout(\processor_zipi8.program_counter_i.un3_half_pcZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNO_1_11_LC_2_13_1 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNO_1_11_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNO_1_11_LC_2_13_1 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNO_1_11_LC_2_13_1  (
            .in0(N__13892),
            .in1(N__21432),
            .in2(N__13883),
            .in3(N__27442),
            .lcout(\processor_zipi8.program_counter_i.un431_half_pc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIKAV8O_2_LC_2_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIKAV8O_2_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNIKAV8O_2_LC_2_13_2 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNIKAV8O_2_LC_2_13_2  (
            .in0(N__15227),
            .in1(N__17773),
            .in2(N__25540),
            .in3(N__17859),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNO_0_11_LC_2_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNO_0_11_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNO_0_11_LC_2_13_4 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNO_0_11_LC_2_13_4  (
            .in0(N__20051),
            .in1(N__14398),
            .in2(N__17871),
            .in3(N__17774),
            .lcout(),
            .ltout(\processor_zipi8.program_counter_i.half_pc_0_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_11_LC_2_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_11_LC_2_13_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_11_LC_2_13_5 .LUT_INIT=16'b1001101011001111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_11_LC_2_13_5  (
            .in0(N__14417),
            .in1(N__14411),
            .in2(N__14405),
            .in3(N__14353),
            .lcout(\processor_zipi8.address_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33635),
            .ce(N__15767),
            .sr(N__17425));
    defparam \processor_zipi8.program_counter_i.pc_RNI70TDO_0_LC_2_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_RNI70TDO_0_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_RNI70TDO_0_LC_2_13_6 .LUT_INIT=16'b0000111011101110;
    LogicCell40 \processor_zipi8.program_counter_i.pc_RNI70TDO_0_LC_2_13_6  (
            .in0(N__15449),
            .in1(N__17772),
            .in2(N__23012),
            .in3(N__17858),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI2ASQ6A_9_LC_2_13_7 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI2ASQ6A_9_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI2ASQ6A_9_LC_2_13_7 .LUT_INIT=16'b1101010100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNI2ASQ6A_9_LC_2_13_7  (
            .in0(N__14387),
            .in1(N__15938),
            .in2(N__14381),
            .in3(N__14365),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_58_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIJJ175_LC_2_14_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIJJ175_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIJJ175_LC_2_14_0 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIJJ175_LC_2_14_0  (
            .in0(N__21179),
            .in1(N__14423),
            .in2(N__18908),
            .in3(N__14432),
            .lcout(\processor_zipi8.pc_mode_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIOK4K1_LC_2_14_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIOK4K1_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIOK4K1_LC_2_14_1 .LUT_INIT=16'b1011011100010010;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIOK4K1_LC_2_14_1  (
            .in0(N__19932),
            .in1(N__14567),
            .in2(N__14342),
            .in3(N__21443),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.N_50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI7M013_LC_2_14_2 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI7M013_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI7M013_LC_2_14_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI7M013_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__14315),
            .in2(N__14333),
            .in3(N__24308),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.N_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIK0IP3_LC_2_14_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIK0IP3_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIK0IP3_LC_2_14_3 .LUT_INIT=16'b0101010111010001;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIK0IP3_LC_2_14_3  (
            .in0(N__14569),
            .in1(N__18874),
            .in2(N__14330),
            .in3(N__21180),
            .lcout(\processor_zipi8.flags_i.N_123_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m44_LC_2_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m44_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m44_LC_2_14_4 .LUT_INIT=16'b0010111110101010;
    LogicCell40 \processor_zipi8.flags_i.m44_LC_2_14_4  (
            .in0(N__21442),
            .in1(N__19931),
            .in2(N__14577),
            .in3(N__24172),
            .lcout(\processor_zipi8.flags_i.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m91_am_LC_2_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m91_am_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m91_am_LC_2_14_5 .LUT_INIT=16'b0110110001100110;
    LogicCell40 \processor_zipi8.flags_i.m91_am_LC_2_14_5  (
            .in0(N__24173),
            .in1(N__14568),
            .in2(N__19958),
            .in3(N__21444),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.m91_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNINARM2_LC_2_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNINARM2_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNINARM2_LC_2_14_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNINARM2_LC_2_14_6  (
            .in0(N__14714),
            .in1(_gnd_net_),
            .in2(N__14441),
            .in3(N__24309),
            .lcout(\processor_zipi8.flags_i.N_1239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m33_LC_2_14_7 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m33_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m33_LC_2_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.flags_i.m33_LC_2_14_7  (
            .in0(N__14491),
            .in1(N__16270),
            .in2(N__14578),
            .in3(N__14657),
            .lcout(\processor_zipi8.flags_i.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNICAJR_0_LC_2_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNICAJR_0_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNICAJR_0_LC_2_15_0 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNICAJR_0_LC_2_15_0  (
            .in0(N__18023),
            .in1(N__24094),
            .in2(_gnd_net_),
            .in3(N__17984),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.m25_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNID1UF1_LC_2_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNID1UF1_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNID1UF1_LC_2_15_1 .LUT_INIT=16'b0011000000000011;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNID1UF1_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__21437),
            .in2(N__14438),
            .in3(N__19901),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.N_26_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI04EE2_LC_2_15_2 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI04EE2_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI04EE2_LC_2_15_2 .LUT_INIT=16'b1111000000010001;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI04EE2_LC_2_15_2  (
            .in0(N__21438),
            .in1(N__24096),
            .in2(N__14435),
            .in3(N__24293),
            .lcout(\processor_zipi8.flags_i.N_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIULO51_LC_2_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIULO51_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIULO51_LC_2_15_3 .LUT_INIT=16'b0001100101011101;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIULO51_LC_2_15_3  (
            .in0(N__24095),
            .in1(N__24291),
            .in2(N__17993),
            .in3(N__18024),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.m20_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIHO842_LC_2_15_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIHO842_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIHO842_LC_2_15_4 .LUT_INIT=16'b1010010111110100;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIHO842_LC_2_15_4  (
            .in0(N__19902),
            .in1(N__21439),
            .in2(N__14426),
            .in3(N__24292),
            .lcout(\processor_zipi8.flags_i.N_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m87_LC_2_15_5 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m87_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m87_LC_2_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \processor_zipi8.flags_i.m87_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__14553),
            .in2(_gnd_net_),
            .in3(N__19903),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.N_1235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI89V91_LC_2_15_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI89V91_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI89V91_LC_2_15_6 .LUT_INIT=16'b0001111011010010;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI89V91_LC_2_15_6  (
            .in0(N__18025),
            .in1(N__24097),
            .in2(N__14717),
            .in3(N__17988),
            .lcout(\processor_zipi8.flags_i.zero_flag_RNI89VZ0Z91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI4LCF3_LC_2_15_7 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI4LCF3_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI4LCF3_LC_2_15_7 .LUT_INIT=16'b0101010111010001;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI4LCF3_LC_2_15_7  (
            .in0(N__14554),
            .in1(N__18913),
            .in2(N__14708),
            .in3(N__21211),
            .lcout(\processor_zipi8.flags_i.N_124_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI281Q3_LC_2_16_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI281Q3_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI281Q3_LC_2_16_0 .LUT_INIT=16'b0011011000000110;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI281Q3_LC_2_16_0  (
            .in0(N__14555),
            .in1(N__16278),
            .in2(N__19069),
            .in3(N__14699),
            .lcout(\processor_zipi8.flags_i.N_1241 ),
            .ltout(\processor_zipi8.flags_i.N_1241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIDS654_LC_2_16_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIDS654_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIDS654_LC_2_16_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIDS654_LC_2_16_1  (
            .in0(N__17402),
            .in1(_gnd_net_),
            .in2(N__14693),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.zero_flag_RNIDS654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.stack_pointer_2_LC_2_16_2 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.stack_pointer_2_LC_2_16_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.stack_pointer_2_LC_2_16_2 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \processor_zipi8.stack_i.stack_pointer_2_LC_2_16_2  (
            .in0(N__19057),
            .in1(N__17405),
            .in2(N__14624),
            .in3(N__14612),
            .lcout(\processor_zipi8.stack_pointer_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33652),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m75_am_LC_2_16_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m75_am_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m75_am_LC_2_16_3 .LUT_INIT=16'b1000000001111111;
    LogicCell40 \processor_zipi8.flags_i.m75_am_LC_2_16_3  (
            .in0(N__16279),
            .in1(N__14662),
            .in2(N__14573),
            .in3(N__14485),
            .lcout(\processor_zipi8.flags_i.m75_amZ0 ),
            .ltout(\processor_zipi8.flags_i.m75_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI5GK75_LC_2_16_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI5GK75_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI5GK75_LC_2_16_4 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI5GK75_LC_2_16_4  (
            .in0(N__19056),
            .in1(N__17403),
            .in2(N__14615),
            .in3(N__14611),
            .lcout(\processor_zipi8.zero_flag_RNI5GK75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.stack_pointer_0_LC_2_16_5 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.stack_pointer_0_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.stack_pointer_0_LC_2_16_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \processor_zipi8.stack_i.stack_pointer_0_LC_2_16_5  (
            .in0(N__17404),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14588),
            .lcout(\processor_zipi8.stack_pointer_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33652),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNI51D94_LC_2_16_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNI51D94_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNI51D94_LC_2_16_6 .LUT_INIT=16'b0101011001000111;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNI51D94_LC_2_16_6  (
            .in0(N__14484),
            .in1(N__16277),
            .in2(N__17259),
            .in3(N__14454),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.m68_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIAKL05_LC_2_16_7 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIAKL05_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIAKL05_LC_2_16_7 .LUT_INIT=16'b1110010010110001;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIAKL05_LC_2_16_7  (
            .in0(N__19009),
            .in1(N__17251),
            .in2(N__14759),
            .in3(N__15102),
            .lcout(\processor_zipi8.flags_i.N_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__6_LC_4_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__6_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__6_LC_4_2_0 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__6_LC_4_2_0  (
            .in0(N__34128),
            .in1(N__36503),
            .in2(N__29329),
            .in3(N__29677),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33654),
            .ce(N__23563),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__7_LC_4_2_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__7_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__7_LC_4_2_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__7_LC_4_2_1  (
            .in0(N__36502),
            .in1(N__33311),
            .in2(N__33009),
            .in3(N__34129),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33654),
            .ce(N__23563),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__6_LC_4_3_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__6_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__6_LC_4_3_0 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__6_LC_4_3_0  (
            .in0(N__34305),
            .in1(N__29201),
            .in2(N__36626),
            .in3(N__29676),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33648),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_6_LC_4_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_6_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_6_LC_4_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_6_LC_4_4_0  (
            .in0(N__16360),
            .in1(N__22376),
            .in2(_gnd_net_),
            .in3(N__37384),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_6_LC_4_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_6_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_6_LC_4_4_1 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_6_LC_4_4_1  (
            .in0(N__14831),
            .in1(N__14735),
            .in2(N__14756),
            .in3(N__28620),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_6_LC_4_4_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_6_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_6_LC_4_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_6_LC_4_4_2  (
            .in0(N__16111),
            .in1(N__16093),
            .in2(_gnd_net_),
            .in3(N__37381),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_6_LC_4_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_6_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_6_LC_4_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_6_LC_4_4_3  (
            .in0(N__37382),
            .in1(N__23809),
            .in2(_gnd_net_),
            .in3(N__16123),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_6_LC_4_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_6_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_6_LC_4_4_4 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_6_LC_4_4_4  (
            .in0(N__28619),
            .in1(N__14744),
            .in2(N__14738),
            .in3(N__29002),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_6_LC_4_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_6_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_6_LC_4_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_6_LC_4_4_5  (
            .in0(N__14921),
            .in1(N__14729),
            .in2(_gnd_net_),
            .in3(N__36034),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268 ),
            .ltout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__6_LC_4_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__6_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__6_LC_4_4_6 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__6_LC_4_4_6  (
            .in0(N__34127),
            .in1(N__29691),
            .in2(N__14834),
            .in3(N__36455),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33644),
            .ce(N__25335),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_6_LC_4_4_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_6_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_6_LC_4_4_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_6_LC_4_4_7  (
            .in0(N__37383),
            .in1(_gnd_net_),
            .in2(N__23462),
            .in3(N__16378),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_0_LC_4_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_0_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_0_LC_4_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_0_LC_4_5_0  (
            .in0(N__14824),
            .in1(N__37078),
            .in2(_gnd_net_),
            .in3(N__14809),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIRJV11_0_LC_4_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIRJV11_0_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIRJV11_0_LC_4_5_1 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIRJV11_0_LC_4_5_1  (
            .in0(N__16510),
            .in1(N__30922),
            .in2(N__31742),
            .in3(N__14792),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIQ8MP1_0_LC_4_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIQ8MP1_0_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIQ8MP1_0_LC_4_5_2 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIQ8MP1_0_LC_4_5_2  (
            .in0(N__14825),
            .in1(N__14810),
            .in2(N__14795),
            .in3(N__31717),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIQ8MP1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_0_LC_4_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_0_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_0_LC_4_5_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_0_LC_4_5_3  (
            .in0(N__37081),
            .in1(_gnd_net_),
            .in2(N__16511),
            .in3(N__14791),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_0_LC_4_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_0_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_0_LC_4_5_4 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_0_LC_4_5_4  (
            .in0(N__28617),
            .in1(N__28978),
            .in2(N__14777),
            .in3(N__14774),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_0_LC_4_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_0_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_0_LC_4_5_5 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_0_LC_4_5_5  (
            .in0(N__14765),
            .in1(N__14882),
            .in2(N__14768),
            .in3(N__28618),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_0_LC_4_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_0_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_0_LC_4_5_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_0_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__18139),
            .in2(N__18121),
            .in3(N__37079),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_0_LC_4_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_0_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_0_LC_4_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_0_LC_4_5_7  (
            .in0(N__37080),
            .in1(N__20387),
            .in2(_gnd_net_),
            .in3(N__20368),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe13_0_a2_LC_4_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe13_0_a2_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe13_0_a2_LC_4_6_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe13_0_a2_LC_4_6_0  (
            .in0(N__20856),
            .in1(N__22246),
            .in2(N__27461),
            .in3(N__20540),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe16_0_a2_LC_4_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe16_0_a2_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe16_0_a2_LC_4_6_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe16_0_a2_LC_4_6_1  (
            .in0(N__27445),
            .in1(N__23153),
            .in2(N__22284),
            .in3(N__20854),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_LC_4_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_LC_4_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_LC_4_6_2  (
            .in0(N__20855),
            .in1(N__22245),
            .in2(N__20326),
            .in3(N__27447),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe8_0_a2_LC_4_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe8_0_a2_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe8_0_a2_LC_4_6_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe8_0_a2_LC_4_6_3  (
            .in0(N__27449),
            .in1(N__23159),
            .in2(N__22287),
            .in3(N__20857),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe10_0_a2_LC_4_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe10_0_a2_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe10_0_a2_LC_4_6_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe10_0_a2_LC_4_6_4  (
            .in0(N__20657),
            .in1(N__22247),
            .in2(N__23163),
            .in3(N__27448),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe18_0_a2_LC_4_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe18_0_a2_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe18_0_a2_LC_4_6_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe18_0_a2_LC_4_6_5  (
            .in0(N__27443),
            .in1(N__23154),
            .in2(N__22286),
            .in3(N__20658),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_LC_4_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_LC_4_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_LC_4_6_6  (
            .in0(N__20659),
            .in1(N__22241),
            .in2(N__23164),
            .in3(N__27446),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe2_0_a2_LC_4_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe2_0_a2_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe2_0_a2_LC_4_6_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe2_0_a2_LC_4_6_7  (
            .in0(N__27444),
            .in1(N__23158),
            .in2(N__22285),
            .in3(N__20660),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe11_0_a2_LC_4_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe11_0_a2_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe11_0_a2_LC_4_7_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe11_0_a2_LC_4_7_0  (
            .in0(N__22138),
            .in1(N__20627),
            .in2(N__20324),
            .in3(N__27455),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe23_0_a2_LC_4_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe23_0_a2_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe23_0_a2_LC_4_7_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe23_0_a2_LC_4_7_1  (
            .in0(N__27451),
            .in1(N__20539),
            .in2(N__20646),
            .in3(N__22135),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe17_0_a2_LC_4_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe17_0_a2_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe17_0_a2_LC_4_7_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe17_0_a2_LC_4_7_2  (
            .in0(N__22134),
            .in1(N__20842),
            .in2(N__20325),
            .in3(N__27453),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe27_0_a2_LC_4_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe27_0_a2_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe27_0_a2_LC_4_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe27_0_a2_LC_4_7_3  (
            .in0(N__27452),
            .in1(N__20316),
            .in2(N__20647),
            .in3(N__22136),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe15_0_a2_LC_4_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe15_0_a2_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe15_0_a2_LC_4_7_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe15_0_a2_LC_4_7_4  (
            .in0(N__22137),
            .in1(N__20628),
            .in2(N__20543),
            .in3(N__27454),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe9_0_a2_LC_4_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe9_0_a2_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe9_0_a2_LC_4_7_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe9_0_a2_LC_4_7_5  (
            .in0(N__27456),
            .in1(N__22139),
            .in2(N__20858),
            .in3(N__20317),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_0_LC_4_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_0_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_0_LC_4_7_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe25_0_a2_0_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__27631),
            .in2(_gnd_net_),
            .in3(N__30984),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212 ),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe1_0_a2_LC_4_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe1_0_a2_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe1_0_a2_LC_4_7_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe1_0_a2_LC_4_7_7  (
            .in0(N__27450),
            .in1(N__20841),
            .in2(N__14885),
            .in3(N__22133),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_0_LC_4_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_0_LC_4_8_0 .SEQ_MODE=4'b1001;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_0_LC_4_8_0 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_0_LC_4_8_0  (
            .in0(N__21702),
            .in1(N__14932),
            .in2(_gnd_net_),
            .in3(N__17129),
            .lcout(\processor_zipi8.shift_rotate_result_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_2_LC_4_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_2_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_2_LC_4_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_2_LC_4_8_1  (
            .in0(N__17128),
            .in1(N__20052),
            .in2(_gnd_net_),
            .in3(N__21701),
            .lcout(\processor_zipi8.shift_rotate_result_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_4_LC_4_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_4_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_4_LC_4_8_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_4_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(N__17127),
            .in2(N__20057),
            .in3(N__18801),
            .lcout(\processor_zipi8.shift_rotate_result_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_6_LC_4_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_6_LC_4_8_3 .SEQ_MODE=4'b1001;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_6_LC_4_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_6_LC_4_8_3  (
            .in0(N__17125),
            .in1(N__16694),
            .in2(_gnd_net_),
            .in3(N__18802),
            .lcout(\processor_zipi8.shift_rotate_result_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_7_LC_4_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_7_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_7_LC_4_8_4 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_7_LC_4_8_4  (
            .in0(N__17124),
            .in1(N__16615),
            .in2(_gnd_net_),
            .in3(N__14933),
            .lcout(\processor_zipi8.shift_rotate_result_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_5_LC_4_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_5_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_5_LC_4_8_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_5_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(N__17122),
            .in2(N__16631),
            .in3(N__21856),
            .lcout(\processor_zipi8.shift_rotate_result_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_3_LC_4_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_3_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_3_LC_4_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_3_LC_4_8_6  (
            .in0(N__21855),
            .in1(N__17126),
            .in2(_gnd_net_),
            .in3(N__22044),
            .lcout(\processor_zipi8.shift_rotate_result_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_1_LC_4_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_1_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_1_LC_4_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_rotate_result_1_LC_4_8_7  (
            .in0(N__22045),
            .in1(N__17123),
            .in2(_gnd_net_),
            .in3(N__21106),
            .lcout(\processor_zipi8.shift_rotate_result_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33612),
            .ce(),
            .sr(N__25796));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_5_0_LC_4_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_5_0_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_5_0_LC_4_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_5_0_LC_4_9_0  (
            .in0(N__14969),
            .in1(N__21441),
            .in2(_gnd_net_),
            .in3(N__25541),
            .lcout(\processor_zipi8.port_id_2 ),
            .ltout(\processor_zipi8.port_id_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_2_LC_4_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_2_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_2_LC_4_9_1 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_2_LC_4_9_1  (
            .in0(N__19577),
            .in1(N__19618),
            .in2(N__14900),
            .in3(N__22040),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_2_LC_4_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_2_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_2_LC_4_9_2 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_2_LC_4_9_2  (
            .in0(N__22041),
            .in1(N__19578),
            .in2(N__15045),
            .in3(N__19180),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_2_LC_4_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_2_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_2_LC_4_9_3 .LUT_INIT=16'b1111111100011011;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_2_LC_4_9_3  (
            .in0(N__15034),
            .in1(N__23999),
            .in2(N__19202),
            .in3(N__22042),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_2_LC_4_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_2_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_2_LC_4_9_4 .LUT_INIT=16'b0001111111111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_2_LC_4_9_4  (
            .in0(N__22039),
            .in1(N__19794),
            .in2(N__19487),
            .in3(N__15035),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_LC_4_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_LC_4_9_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_LC_4_9_5  (
            .in0(N__15011),
            .in1(N__15005),
            .in2(N__14999),
            .in3(N__14996),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI9VF21_2_LC_4_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI9VF21_2_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI9VF21_2_LC_4_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI9VF21_2_LC_4_9_6  (
            .in0(N__14990),
            .in1(N__14968),
            .in2(_gnd_net_),
            .in3(N__21440),
            .lcout(\processor_zipi8.pc_vector_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_RNO_5_LC_4_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_5_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_5_LC_4_9_7 .LUT_INIT=16'b0110100110100101;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_RNO_5_LC_4_9_7  (
            .in0(N__32324),
            .in1(N__21227),
            .in2(N__39546),
            .in3(N__17990),
            .lcout(\processor_zipi8.flags_i.parity_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_3_LC_4_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_3_LC_4_10_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_3_LC_4_10_0 .LUT_INIT=16'b0000001011111101;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_3_LC_4_10_0  (
            .in0(N__15350),
            .in1(N__15371),
            .in2(N__15980),
            .in3(N__15869),
            .lcout(address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33630),
            .ce(N__15758),
            .sr(N__17390));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_LC_4_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_LC_4_10_1 .LUT_INIT=16'b0011110111111101;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_LC_4_10_1  (
            .in0(N__17991),
            .in1(N__21516),
            .in2(N__14975),
            .in3(N__17002),
            .lcout(),
            .ltout(\processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_1_LC_4_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_1_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_1_LC_4_10_2 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_1_LC_4_10_2  (
            .in0(N__21517),
            .in1(N__16702),
            .in2(N__14978),
            .in3(N__14973),
            .lcout(),
            .ltout(\processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_LC_4_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_LC_4_10_3 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \processor_zipi8.shift_and_rotate_operations_i.shift_in_bit_LC_4_10_3  (
            .in0(N__14974),
            .in1(N__21518),
            .in2(N__14936),
            .in3(N__21090),
            .lcout(\processor_zipi8.shift_and_rotate_operations_i.shift_in_bitZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_1_LC_4_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_1_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_1_LC_4_10_4 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \processor_zipi8.register_bank_control_i.bank_RNO_1_LC_4_10_4  (
            .in0(N__16049),
            .in1(N__17543),
            .in2(N__19059),
            .in3(N__16718),
            .lcout(\processor_zipi8.register_bank_control_i.un1_bank_value ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_2_LC_4_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_2_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_esr_2_LC_4_10_5 .LUT_INIT=16'b0110011000110011;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_2_LC_4_10_5  (
            .in0(N__15370),
            .in1(N__15976),
            .in2(_gnd_net_),
            .in3(N__15349),
            .lcout(address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33630),
            .ce(N__15758),
            .sr(N__17390));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5LPHH_0_LC_4_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5LPHH_0_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5LPHH_0_LC_4_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5LPHH_0_LC_4_10_6  (
            .in0(N__22132),
            .in1(N__24779),
            .in2(_gnd_net_),
            .in3(N__20555),
            .lcout(\processor_zipi8.sx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m57_LC_4_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m57_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m57_LC_4_11_0 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \processor_zipi8.flags_i.m57_LC_4_11_0  (
            .in0(N__17230),
            .in1(N__15157),
            .in2(_gnd_net_),
            .in3(N__15109),
            .lcout(\processor_zipi8.flags_i.i14_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_RNO_0_0_LC_4_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_RNO_0_0_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_RNO_0_0_LC_4_11_1 .LUT_INIT=16'b0111101100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_RNO_0_0_LC_4_11_1  (
            .in0(N__16013),
            .in1(N__15956),
            .in2(N__15062),
            .in3(N__15842),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_7_0_LC_4_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_7_0_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_7_0_LC_4_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_7_0_LC_4_11_2  (
            .in0(N__21401),
            .in1(N__17000),
            .in2(_gnd_net_),
            .in3(N__23005),
            .lcout(\processor_zipi8.port_id_0 ),
            .ltout(\processor_zipi8.port_id_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_LC_4_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_LC_4_11_3 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_LC_4_11_3  (
            .in0(N__19457),
            .in1(N__19783),
            .in2(N__15083),
            .in3(N__21083),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_1_LC_4_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_1_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_1_LC_4_11_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_1_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__17030),
            .in2(_gnd_net_),
            .in3(N__19283),
            .lcout(\processor_zipi8.arith_logical_result_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33637),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_0_LC_4_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_0_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_0_LC_4_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_0_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15080),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33637),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI6TF21_0_LC_4_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI6TF21_0_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI6TF21_0_LC_4_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI6TF21_0_LC_4_11_6  (
            .in0(N__21402),
            .in1(N__15068),
            .in2(_gnd_net_),
            .in3(N__17001),
            .lcout(\processor_zipi8.pc_vector_0 ),
            .ltout(\processor_zipi8.pc_vector_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_RNIUJNL41_0_LC_4_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_RNIUJNL41_0_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_RNIUJNL41_0_LC_4_11_7 .LUT_INIT=16'b0101000100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_RNIUJNL41_0_LC_4_11_7  (
            .in0(N__16012),
            .in1(N__15955),
            .in2(N__15845),
            .in3(N__15841),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNIC4FP9_LC_4_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIC4FP9_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIC4FP9_LC_4_12_0 .LUT_INIT=16'b0000000101000101;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIC4FP9_LC_4_12_0  (
            .in0(N__17414),
            .in1(N__19066),
            .in2(N__15826),
            .in3(N__15802),
            .lcout(\processor_zipi8.zero_flag_RNIC4FP9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_ctle_11_LC_4_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_ctle_11_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_ctle_11_LC_4_12_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_ctle_11_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__17412),
            .in2(_gnd_net_),
            .in3(N__19065),
            .lcout(\processor_zipi8.program_counter_i.t_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_RNI72UDO_1_LC_4_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_RNI72UDO_1_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_RNI72UDO_1_LC_4_12_2 .LUT_INIT=16'b0100010111001111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_RNI72UDO_1_LC_4_12_2  (
            .in0(N__17850),
            .in1(N__17798),
            .in2(N__15611),
            .in3(N__23198),
            .lcout(),
            .ltout(\processor_zipi8.program_counter_i.half_pc_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_RNINDAA01_1_LC_4_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_RNINDAA01_1_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_RNINDAA01_1_LC_4_12_3 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_RNINDAA01_1_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__21482),
            .in2(N__15722),
            .in3(N__15957),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_1 ),
            .ltout(\processor_zipi8.program_counter_i.half_pc_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_1_LC_4_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_1_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_1_LC_4_12_4 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \processor_zipi8.program_counter_i.pc_1_LC_4_12_4  (
            .in0(N__15348),
            .in1(N__15602),
            .in2(N__15719),
            .in3(N__19068),
            .lcout(address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33643),
            .ce(),
            .sr(N__17415));
    defparam \processor_zipi8.program_counter_i.pc_0_LC_4_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_0_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.program_counter_i.pc_0_LC_4_12_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \processor_zipi8.program_counter_i.pc_0_LC_4_12_5  (
            .in0(N__19067),
            .in1(N__15548),
            .in2(_gnd_net_),
            .in3(N__15441),
            .lcout(address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33643),
            .ce(),
            .sr(N__17415));
    defparam \processor_zipi8.flags_i.zero_flag_RNIL8RB5_LC_4_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNIL8RB5_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNIL8RB5_LC_4_12_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNIL8RB5_LC_4_12_6  (
            .in0(N__17413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17281),
            .lcout(\processor_zipi8.zero_flag_RNIL8RB5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI3JQA54_3_LC_4_12_7 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI3JQA54_3_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI3JQA54_3_LC_4_12_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNI3JQA54_3_LC_4_12_7  (
            .in0(N__15970),
            .in1(N__15865),
            .in2(N__15369),
            .in3(N__15347),
            .lcout(\processor_zipi8.program_counter_i.carry_pc_22_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_LC_4_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_LC_4_13_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_LC_4_13_0  (
            .in0(N__24153),
            .in1(N__16730),
            .in2(N__18883),
            .in3(N__24276),
            .lcout(\processor_zipi8.pc_mode_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI6NB501_2_LC_4_13_1 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI6NB501_2_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI6NB501_2_LC_4_13_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNI6NB501_2_LC_4_13_1  (
            .in0(N__15998),
            .in1(N__15958),
            .in2(_gnd_net_),
            .in3(N__15989),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8QC501_3_LC_4_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8QC501_3_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNI8QC501_3_LC_4_13_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNI8QC501_3_LC_4_13_2  (
            .in0(N__15959),
            .in1(N__17054),
            .in2(_gnd_net_),
            .in3(N__17573),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_1_LC_4_13_3 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_1_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_1_LC_4_13_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \processor_zipi8.decode4alu_i.arith_logical_sel_1_1_LC_4_13_3  (
            .in0(N__24275),
            .in1(N__19944),
            .in2(_gnd_net_),
            .in3(N__24154),
            .lcout(\processor_zipi8.arith_logical_sel_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m101_e_LC_4_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m101_e_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m101_e_LC_4_13_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \processor_zipi8.flags_i.m101_e_LC_4_13_4  (
            .in0(N__24155),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24277),
            .lcout(\processor_zipi8.un16_alu_mux_sel_value ),
            .ltout(\processor_zipi8.un16_alu_mux_sel_value_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.register_bank_control_i.sx_addr_4_LC_4_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.register_bank_control_i.sx_addr_4_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.register_bank_control_i.sx_addr_4_LC_4_13_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \processor_zipi8.register_bank_control_i.sx_addr_4_LC_4_13_5  (
            .in0(N__16133),
            .in1(_gnd_net_),
            .in2(N__15854),
            .in3(N__25609),
            .lcout(\processor_zipi8.sx_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33647),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_4_LC_4_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_4_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_4_LC_4_13_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_4_LC_4_13_6  (
            .in0(N__21216),
            .in1(N__24161),
            .in2(N__18884),
            .in3(N__24278),
            .lcout(\processor_zipi8.decode4_strobes_enables_i.un23_flag_enable_type ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_pc_statck_i.returni_type_o_2_LC_4_13_7 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_pc_statck_i.returni_type_o_2_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_pc_statck_i.returni_type_o_2_LC_4_13_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \processor_zipi8.decode4_pc_statck_i.returni_type_o_2_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__21215),
            .in2(_gnd_net_),
            .in3(N__19945),
            .lcout(\processor_zipi8.returni_type_o_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_3_LC_4_14_0 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_3_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_3_LC_4_14_0 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_3_LC_4_14_0  (
            .in0(N__21224),
            .in1(N__19937),
            .in2(N__18931),
            .in3(N__15851),
            .lcout(),
            .ltout(\processor_zipi8.decode4_strobes_enables_i.flag_enable_type_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_1_LC_4_14_1 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_1_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_1_LC_4_14_1 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_1_LC_4_14_1  (
            .in0(N__19938),
            .in1(N__18921),
            .in2(N__16076),
            .in3(N__24289),
            .lcout(\processor_zipi8.decode4_strobes_enables_i.flag_enable_type_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_2_LC_4_14_2 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_2_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_2_LC_4_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_2_LC_4_14_2  (
            .in0(N__16073),
            .in1(N__16064),
            .in2(_gnd_net_),
            .in3(N__35731),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_4_LC_4_14_3 .C_ON=1'b0;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_4_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_4_LC_4_14_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.register_bank_control_i.bank_RNO_4_LC_4_14_3  (
            .in0(N__19936),
            .in1(N__21223),
            .in2(N__21457),
            .in3(N__24288),
            .lcout(),
            .ltout(\processor_zipi8.register_bank_control_i.un31_regbank_type_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_3_LC_4_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_3_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_3_LC_4_14_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \processor_zipi8.register_bank_control_i.bank_RNO_3_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__18914),
            .in2(N__16052),
            .in3(N__24170),
            .lcout(\processor_zipi8.register_bank_control_i.un31_regbank_type ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.spm_enable_RNO_0_LC_4_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.spm_enable_RNO_0_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.spm_enable_RNO_0_LC_4_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.spm_enable_RNO_0_LC_4_14_5  (
            .in0(N__19939),
            .in1(N__21225),
            .in2(N__18930),
            .in3(N__19060),
            .lcout(\processor_zipi8.decode4_strobes_enables_i.spm_enable_value_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_0_LC_4_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_0_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_0_LC_4_14_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_0_LC_4_14_6  (
            .in0(N__16040),
            .in1(N__35730),
            .in2(_gnd_net_),
            .in3(N__16031),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_1_LC_4_14_7 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_1_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_1_LC_4_14_7 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \processor_zipi8.decode4alu_i.alu_mux_sel_1_LC_4_14_7  (
            .in0(N__24171),
            .in1(_gnd_net_),
            .in2(N__19959),
            .in3(N__24290),
            .lcout(\processor_zipi8.alu_mux_sel_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33653),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_LC_4_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_LC_4_15_0 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_LC_4_15_0  (
            .in0(N__16304),
            .in1(N__17924),
            .in2(N__18929),
            .in3(N__24331),
            .lcout(),
            .ltout(\processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_LC_4_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_LC_4_15_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \processor_zipi8.decode4_pc_statck_i.pc_mode_2_0_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16016),
            .in3(N__16298),
            .lcout(\processor_zipi8.pc_mode_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_pc_statck_i.un3_pc_mode_LC_4_15_2 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_pc_statck_i.un3_pc_mode_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_pc_statck_i.un3_pc_mode_LC_4_15_2 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \processor_zipi8.decode4_pc_statck_i.un3_pc_mode_LC_4_15_2  (
            .in0(N__21416),
            .in1(N__24327),
            .in2(N__24169),
            .in3(N__21181),
            .lcout(\processor_zipi8.decode4_pc_statck_i.un3_pc_modeZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m16_LC_4_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m16_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m16_LC_4_15_3 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \processor_zipi8.flags_i.m16_LC_4_15_3  (
            .in0(N__24147),
            .in1(N__21417),
            .in2(N__24340),
            .in3(N__19946),
            .lcout(\processor_zipi8.N_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.m104_2_LC_4_15_5 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.m104_2_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.m104_2_LC_4_15_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \processor_zipi8.flags_i.m104_2_LC_4_15_5  (
            .in0(N__21182),
            .in1(N__18912),
            .in2(N__16292),
            .in3(N__19947),
            .lcout(\processor_zipi8.flags_i.m104Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__7_LC_5_1_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__7_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__7_LC_5_1_0 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__7_LC_5_1_0  (
            .in0(N__36688),
            .in1(N__34571),
            .in2(N__33342),
            .in3(N__33016),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33668),
            .ce(N__24917),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__6_LC_5_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__6_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__6_LC_5_2_0 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__6_LC_5_2_0  (
            .in0(N__34130),
            .in1(N__36484),
            .in2(N__29367),
            .in3(N__29675),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33662),
            .ce(N__20141),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__7_LC_5_2_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__7_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__7_LC_5_2_1 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__7_LC_5_2_1  (
            .in0(N__34569),
            .in1(N__33309),
            .in2(N__33014),
            .in3(N__36501),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33662),
            .ce(N__20141),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__4_LC_5_3_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__4_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__4_LC_5_3_7 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__4_LC_5_3_7  (
            .in0(N__34306),
            .in1(N__35193),
            .in2(N__36848),
            .in3(N__35427),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33655),
            .ce(N__32674),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNINVTE1_6_LC_5_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNINVTE1_6_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNINVTE1_6_LC_5_4_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNINVTE1_6_LC_5_4_0  (
            .in0(N__16124),
            .in1(N__31590),
            .in2(N__23813),
            .in3(N__30932),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI44F42_6_LC_5_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI44F42_6_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI44F42_6_LC_5_4_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI44F42_6_LC_5_4_1  (
            .in0(N__31591),
            .in1(N__16112),
            .in2(N__16100),
            .in3(N__16097),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNI44F42_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMVAG4_6_LC_5_4_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMVAG4_6_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMVAG4_6_LC_5_4_2 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMVAG4_6_LC_5_4_2  (
            .in0(N__27386),
            .in1(N__16343),
            .in2(N__16079),
            .in3(N__27640),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIVVE01_6_LC_5_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIVVE01_6_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIVVE01_6_LC_5_4_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIVVE01_6_LC_5_4_3  (
            .in0(N__30931),
            .in1(N__23461),
            .in2(N__31695),
            .in3(N__16379),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIK4HN1_6_LC_5_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIK4HN1_6_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIK4HN1_6_LC_5_4_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIK4HN1_6_LC_5_4_4  (
            .in0(N__22375),
            .in1(N__16361),
            .in2(N__16346),
            .in3(N__31589),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIK4HN1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7B4G8_6_LC_5_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7B4G8_6_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7B4G8_6_LC_5_4_5 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7B4G8_6_LC_5_4_5  (
            .in0(N__16337),
            .in1(N__16328),
            .in2(N__16322),
            .in3(N__27387),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7B4G8_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5RVHH_6_LC_5_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5RVHH_6_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5RVHH_6_LC_5_4_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5RVHH_6_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__22415),
            .in2(N__16307),
            .in3(N__22234),
            .lcout(\processor_zipi8.sx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__0_LC_5_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__0_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__0_LC_5_5_0 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__0_LC_5_5_0  (
            .in0(N__36705),
            .in1(N__33951),
            .in2(N__32098),
            .in3(N__32240),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__1_LC_5_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__1_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__1_LC_5_5_1 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__1_LC_5_5_1  (
            .in0(N__33947),
            .in1(N__36709),
            .in2(N__39262),
            .in3(N__39591),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__2_LC_5_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__2_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__2_LC_5_5_2 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__2_LC_5_5_2  (
            .in0(N__36706),
            .in1(N__33952),
            .in2(N__38881),
            .in3(N__38462),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__3_LC_5_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__3_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__3_LC_5_5_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__3_LC_5_5_3  (
            .in0(N__33948),
            .in1(N__36710),
            .in2(N__37824),
            .in3(N__38098),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__4_LC_5_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__4_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__4_LC_5_5_4 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__4_LC_5_5_4  (
            .in0(N__36707),
            .in1(N__33954),
            .in2(N__35191),
            .in3(N__35549),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__5_LC_5_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__5_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__5_LC_5_5_5 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__5_LC_5_5_5  (
            .in0(N__33949),
            .in1(N__36711),
            .in2(N__30463),
            .in3(N__30076),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__6_LC_5_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__6_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__6_LC_5_5_6 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__6_LC_5_5_6  (
            .in0(N__36708),
            .in1(N__33953),
            .in2(N__29704),
            .in3(N__29357),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__7_LC_5_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__7_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__7_LC_5_5_7 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram13__7_LC_5_5_7  (
            .in0(N__33950),
            .in1(N__36712),
            .in2(N__32994),
            .in3(N__33256),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33645),
            .ce(N__16409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__0_LC_5_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__0_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__0_LC_5_6_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__0_LC_5_6_0  (
            .in0(N__34499),
            .in1(N__32380),
            .in2(N__32097),
            .in3(N__36814),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__1_LC_5_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__1_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__1_LC_5_6_1 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__1_LC_5_6_1  (
            .in0(N__36807),
            .in1(N__39247),
            .in2(N__39593),
            .in3(N__34505),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__2_LC_5_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__2_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__2_LC_5_6_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__2_LC_5_6_2  (
            .in0(N__34500),
            .in1(N__36811),
            .in2(N__38532),
            .in3(N__38886),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__3_LC_5_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__3_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__3_LC_5_6_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__3_LC_5_6_3  (
            .in0(N__36808),
            .in1(N__34503),
            .in2(N__38158),
            .in3(N__37701),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__4_LC_5_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__4_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__4_LC_5_6_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__4_LC_5_6_4  (
            .in0(N__34501),
            .in1(N__36812),
            .in2(N__35192),
            .in3(N__35426),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__5_LC_5_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__5_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__5_LC_5_6_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__5_LC_5_6_5  (
            .in0(N__36809),
            .in1(N__30386),
            .in2(N__30137),
            .in3(N__34506),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__6_LC_5_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__6_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__6_LC_5_6_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__6_LC_5_6_6  (
            .in0(N__34502),
            .in1(N__36813),
            .in2(N__29301),
            .in3(N__29554),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__7_LC_5_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__7_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__7_LC_5_6_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__7_LC_5_6_7  (
            .in0(N__36810),
            .in1(N__33266),
            .in2(N__33012),
            .in3(N__34504),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33638),
            .ce(N__16523),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__0_LC_5_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__0_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__0_LC_5_7_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__0_LC_5_7_0  (
            .in0(N__34507),
            .in1(N__32244),
            .in2(N__32099),
            .in3(N__36699),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__1_LC_5_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__1_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__1_LC_5_7_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__1_LC_5_7_1  (
            .in0(N__36692),
            .in1(N__34511),
            .in2(N__39597),
            .in3(N__39094),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__2_LC_5_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__2_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__2_LC_5_7_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__2_LC_5_7_2  (
            .in0(N__34508),
            .in1(N__36698),
            .in2(N__38540),
            .in3(N__38851),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__3_LC_5_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__3_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__3_LC_5_7_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__3_LC_5_7_3  (
            .in0(N__36693),
            .in1(N__38099),
            .in2(N__37853),
            .in3(N__34512),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__4_LC_5_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__4_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__4_LC_5_7_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__4_LC_5_7_4  (
            .in0(N__34509),
            .in1(N__36696),
            .in2(N__35218),
            .in3(N__35511),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__5_LC_5_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__5_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__5_LC_5_7_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__5_LC_5_7_5  (
            .in0(N__36694),
            .in1(N__30394),
            .in2(N__30044),
            .in3(N__34513),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__6_LC_5_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__6_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__6_LC_5_7_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__6_LC_5_7_6  (
            .in0(N__34510),
            .in1(N__36697),
            .in2(N__29364),
            .in3(N__29553),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__7_LC_5_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__7_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__7_LC_5_7_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__7_LC_5_7_7  (
            .in0(N__36695),
            .in1(N__33174),
            .in2(N__33029),
            .in3(N__34514),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33631),
            .ce(N__16454),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__0_LC_5_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__0_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__0_LC_5_8_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__0_LC_5_8_0  (
            .in0(N__34516),
            .in1(N__36413),
            .in2(N__32299),
            .in3(N__31988),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33621),
            .ce(N__18083),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__1_LC_5_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__1_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__1_LC_5_8_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__1_LC_5_8_1  (
            .in0(N__36410),
            .in1(N__34518),
            .in2(N__39594),
            .in3(N__39052),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33621),
            .ce(N__18083),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__2_LC_5_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__2_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__2_LC_5_8_2 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__2_LC_5_8_2  (
            .in0(N__38545),
            .in1(N__36414),
            .in2(N__38880),
            .in3(N__34515),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33621),
            .ce(N__18083),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__3_LC_5_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__3_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__3_LC_5_8_3 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__3_LC_5_8_3  (
            .in0(N__36411),
            .in1(N__38123),
            .in2(N__34700),
            .in3(N__37801),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33621),
            .ce(N__18083),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__4_LC_5_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__4_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__4_LC_5_8_4 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__4_LC_5_8_4  (
            .in0(N__34517),
            .in1(N__35363),
            .in2(N__36607),
            .in3(N__35006),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33621),
            .ce(N__18083),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__5_LC_5_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__5_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__5_LC_5_8_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__5_LC_5_8_5  (
            .in0(N__36412),
            .in1(N__34519),
            .in2(N__30462),
            .in3(N__30057),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33621),
            .ce(N__18083),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_3_0_LC_5_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_3_0_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_3_0_LC_5_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_3_0_LC_5_8_7  (
            .in0(N__16949),
            .in1(N__21445),
            .in2(_gnd_net_),
            .in3(N__37486),
            .lcout(\processor_zipi8.port_id_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.arith_carry_LC_5_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.arith_carry_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.flags_i.arith_carry_LC_5_9_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \processor_zipi8.flags_i.arith_carry_LC_5_9_0  (
            .in0(N__19796),
            .in1(N__16553),
            .in2(N__16706),
            .in3(N__16562),
            .lcout(\processor_zipi8.flags_i.arith_carryZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33632),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical6_process_carry_arith_logical_40_6_LC_5_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical6_process_carry_arith_logical_40_6_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical6_process_carry_arith_logical_40_6_LC_5_9_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical6_process_carry_arith_logical_40_6_LC_5_9_1  (
            .in0(N__16798),
            .in1(N__19795),
            .in2(N__16619),
            .in3(N__19330),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6 ),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_40_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_7_LC_5_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_7_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_7_LC_5_9_2 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_7_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16556),
            .in3(N__16552),
            .lcout(\processor_zipi8.arith_logical_result_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33632),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_6_LC_5_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_6_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_6_LC_5_9_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_6_LC_5_9_3  (
            .in0(N__16799),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19331),
            .lcout(\processor_zipi8.arith_logical_result_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33632),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_RNO_3_LC_5_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_3_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_3_LC_5_9_4 .LUT_INIT=16'b0011011111110111;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_RNO_3_LC_5_9_4  (
            .in0(N__16769),
            .in1(N__16910),
            .in2(N__19964),
            .in3(N__16756),
            .lcout(),
            .ltout(\processor_zipi8.flags_i.carry_flag_value_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_RNO_0_LC_5_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_0_LC_5_9_5 .LUT_INIT=16'b1101000000000000;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_RNO_0_LC_5_9_5  (
            .in0(N__16712),
            .in1(N__16775),
            .in2(N__16784),
            .in3(N__16736),
            .lcout(\processor_zipi8.flags_i.carry_flag_value_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_RNO_1_LC_5_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_1_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_1_LC_5_9_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_RNO_1_LC_5_9_6  (
            .in0(N__29499),
            .in1(N__19304),
            .in2(N__33147),
            .in3(N__16781),
            .lcout(\processor_zipi8.flags_i.carry_flag_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_RNO_2_LC_5_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_2_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_2_LC_5_9_7 .LUT_INIT=16'b0010101000111111;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_RNO_2_LC_5_9_7  (
            .in0(N__16768),
            .in1(N__16879),
            .in2(N__16757),
            .in3(N__23986),
            .lcout(\processor_zipi8.flags_i.carry_flag_value_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un52_half_arith_logical_LC_5_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un52_half_arith_logical_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un52_half_arith_logical_LC_5_10_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un52_half_arith_logical_LC_5_10_0  (
            .in0(N__19779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19186),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.un52_half_arith_logical ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_1_LC_5_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_1_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_1_LC_5_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \processor_zipi8.decode4_pc_statck_i.un47_pc_mode_1_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__21399),
            .in2(_gnd_net_),
            .in3(N__19949),
            .lcout(\processor_zipi8.decode4_pc_statck_i.N_22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_2_LC_5_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_2_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_2_LC_5_10_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.register_bank_control_i.bank_RNO_2_LC_5_10_2  (
            .in0(N__21400),
            .in1(N__24323),
            .in2(N__18932),
            .in3(N__24163),
            .lcout(\processor_zipi8.register_bank_control_i.un17_regbank_type_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_RNO_4_LC_5_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_4_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_4_LC_5_10_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_RNO_4_LC_5_10_3  (
            .in0(N__24164),
            .in1(_gnd_net_),
            .in2(N__24338),
            .in3(N__19951),
            .lcout(\processor_zipi8.flags_i.un17_carry_flag_value_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_value_1_LC_5_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_value_1_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_value_1_LC_5_10_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \processor_zipi8.decode4alu_i.alu_mux_sel_value_1_LC_5_10_4  (
            .in0(N__19950),
            .in1(N__24319),
            .in2(_gnd_net_),
            .in3(N__24162),
            .lcout(\processor_zipi8.alu_mux_sel_value_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_1_LC_5_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_1_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_1_LC_5_10_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_1_LC_5_10_5  (
            .in0(N__24165),
            .in1(_gnd_net_),
            .in2(N__24339),
            .in3(N__17542),
            .lcout(\processor_zipi8.decode4_strobes_enables_i.un8_register_enable_type ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical2_process_carry_arith_logical_16_2_LC_5_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical2_process_carry_arith_logical_16_2_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical2_process_carry_arith_logical_16_2_LC_5_10_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical2_process_carry_arith_logical_16_2_LC_5_10_6  (
            .in0(N__19780),
            .in1(N__16861),
            .in2(N__22043),
            .in3(N__17014),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2 ),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_16_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical3_process_carry_arith_logical_22_3_LC_5_10_7 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical3_process_carry_arith_logical_22_3_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical3_process_carry_arith_logical_22_3_LC_5_10_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical3_process_carry_arith_logical_22_3_LC_5_10_7  (
            .in0(N__20050),
            .in1(N__19102),
            .in2(N__16850),
            .in3(N__19781),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_22_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_21_tz_LC_5_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_21_tz_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_21_tz_LC_5_11_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_21_tz_LC_5_11_0  (
            .in0(N__19467),
            .in1(N__19187),
            .in2(_gnd_net_),
            .in3(N__21685),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.N_773_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_0_LC_5_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_0_LC_5_11_1 .LUT_INIT=16'b1001110111111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_0_LC_5_11_1  (
            .in0(N__19188),
            .in1(N__21078),
            .in2(N__19778),
            .in3(N__16821),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_0_LC_5_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_0_LC_5_11_2 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_0_LC_5_11_2  (
            .in0(N__21079),
            .in1(N__16823),
            .in2(N__16847),
            .in3(N__23988),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_0_LC_5_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_0_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_0_LC_5_11_3 .LUT_INIT=16'b1101000001110000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_0_LC_5_11_3  (
            .in0(N__19557),
            .in1(N__21080),
            .in2(N__16844),
            .in3(N__16822),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un36_half_arith_logical_1_LC_5_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un36_half_arith_logical_1_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un36_half_arith_logical_1_LC_5_11_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_half_arith_logical0_process_un36_half_arith_logical_1_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__16824),
            .in2(_gnd_net_),
            .in3(N__19189),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.un36_half_arith_logical_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_LC_5_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_LC_5_11_5 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_LC_5_11_5  (
            .in0(N__19294),
            .in1(N__21081),
            .in2(N__17048),
            .in3(N__17039),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0 ),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical0_process_carry_arith_logical_4_0_LC_5_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical0_process_carry_arith_logical_4_0_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical0_process_carry_arith_logical_4_0_LC_5_11_6 .LUT_INIT=16'b0000001110100011;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical0_process_carry_arith_logical_4_0_LC_5_11_6  (
            .in0(N__21082),
            .in1(N__17563),
            .in2(N__17033),
            .in3(N__19743),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0 ),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical1_process_carry_arith_logical_10_1_LC_5_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical1_process_carry_arith_logical_10_1_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical1_process_carry_arith_logical_10_1_LC_5_11_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical1_process_carry_arith_logical_10_1_LC_5_11_7  (
            .in0(N__21686),
            .in1(N__19784),
            .in2(N__17024),
            .in3(N__19279),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_0_LC_5_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_0_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.register_bank_control_i.bank_RNO_0_LC_5_12_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \processor_zipi8.register_bank_control_i.bank_RNO_0_LC_5_12_0  (
            .in0(N__24314),
            .in1(N__16916),
            .in2(_gnd_net_),
            .in3(N__17003),
            .lcout(),
            .ltout(\processor_zipi8.register_bank_control_i.bank_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.register_bank_control_i.bank_LC_5_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.register_bank_control_i.bank_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.register_bank_control_i.bank_LC_5_12_1 .LUT_INIT=16'b1010101000101110;
    LogicCell40 \processor_zipi8.register_bank_control_i.bank_LC_5_12_1  (
            .in0(N__25605),
            .in1(N__16964),
            .in2(N__16952),
            .in3(N__17442),
            .lcout(\processor_zipi8.bank ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33649),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_4_LC_5_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_4_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_4_LC_5_12_2 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_4_LC_5_12_2  (
            .in0(N__19343),
            .in1(N__19970),
            .in2(N__24590),
            .in3(N__25604),
            .lcout(\processor_zipi8.sy_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.shadow_carry_flag_2_LC_5_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_2_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.shadow_carry_flag_2_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \processor_zipi8.stack_i.shadow_carry_flag_2_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16931),
            .lcout(\processor_zipi8.shadow_bank ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33649),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.calc_arith_logical_sel_process_un4_arith_logical_sel_LC_5_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.calc_arith_logical_sel_process_un4_arith_logical_sel_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4alu_i.calc_arith_logical_sel_process_un4_arith_logical_sel_LC_5_12_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \processor_zipi8.decode4alu_i.calc_arith_logical_sel_process_un4_arith_logical_sel_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__16903),
            .in2(_gnd_net_),
            .in3(N__19948),
            .lcout(\processor_zipi8.un4_arith_logical_sel ),
            .ltout(\processor_zipi8.un4_arith_logical_sel_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.arith_carry_in_LC_5_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.arith_carry_in_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4alu_i.arith_carry_in_LC_5_12_5 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \processor_zipi8.decode4alu_i.arith_carry_in_LC_5_12_5  (
            .in0(N__21214),
            .in1(N__23976),
            .in2(N__16892),
            .in3(N__17959),
            .lcout(\processor_zipi8.arith_carry_in_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_LC_5_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.flags_i.carry_flag_LC_5_12_6 .LUT_INIT=16'b0000001000110010;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_LC_5_12_6  (
            .in0(N__17960),
            .in1(N__17443),
            .in2(N__17507),
            .in3(N__17453),
            .lcout(\processor_zipi8.carry_flag ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33649),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.stack_i.stack_pointer_3_LC_5_12_7 .C_ON=1'b0;
    defparam \processor_zipi8.stack_i.stack_pointer_3_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.stack_i.stack_pointer_3_LC_5_12_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \processor_zipi8.stack_i.stack_pointer_3_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__17441),
            .in2(_gnd_net_),
            .in3(N__17285),
            .lcout(\processor_zipi8.stack_pointer_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33649),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_3_LC_5_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_3_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_3_LC_5_13_0 .LUT_INIT=16'b0101001111111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0_3_LC_5_13_0  (
            .in0(N__19631),
            .in1(N__19551),
            .in2(N__20046),
            .in3(N__17156),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_LC_5_13_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_LC_5_13_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_LC_5_13_1  (
            .in0(N__17135),
            .in1(N__17201),
            .in2(N__17204),
            .in3(N__17192),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_3_LC_5_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_3_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_3_LC_5_13_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_3_LC_5_13_2  (
            .in0(N__19563),
            .in1(N__17155),
            .in2(N__20045),
            .in3(N__19153),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_4_0_LC_5_13_3 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_4_0_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_4_0_LC_5_13_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_4_0_LC_5_13_3  (
            .in0(N__17101),
            .in1(N__21356),
            .in2(_gnd_net_),
            .in3(N__19652),
            .lcout(\processor_zipi8.port_id_3 ),
            .ltout(\processor_zipi8.port_id_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_3_LC_5_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_3_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_3_LC_5_13_4 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_3_LC_5_13_4  (
            .in0(N__19473),
            .in1(N__20014),
            .in2(N__17195),
            .in3(N__19739),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_3_LC_5_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_3_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_3_LC_5_13_5 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2_3_LC_5_13_5  (
            .in0(N__19152),
            .in1(N__20024),
            .in2(N__17166),
            .in3(N__23985),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIA0G21_3_LC_5_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIA0G21_3_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIA0G21_3_LC_5_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIA0G21_3_LC_5_13_6  (
            .in0(N__21355),
            .in1(N__23633),
            .in2(_gnd_net_),
            .in3(N__17100),
            .lcout(\processor_zipi8.pc_vector_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.program_counter_i.pc_esr_RNILC09O_3_LC_5_13_7 .C_ON=1'b0;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNILC09O_3_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.program_counter_i.pc_esr_RNILC09O_3_LC_5_13_7 .LUT_INIT=16'b0100010111001111;
    LogicCell40 \processor_zipi8.program_counter_i.pc_esr_RNILC09O_3_LC_5_13_7  (
            .in0(N__17849),
            .in1(N__17804),
            .in2(N__17640),
            .in3(N__19651),
            .lcout(\processor_zipi8.program_counter_i.half_pc_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_0_LC_5_14_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_0_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_0_LC_5_14_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_0_LC_5_14_2  (
            .in0(N__17567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17552),
            .lcout(\processor_zipi8.arith_logical_result_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33661),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_2_LC_5_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_2_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_2_LC_5_14_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_2_LC_5_14_4  (
            .in0(N__17530),
            .in1(N__18927),
            .in2(_gnd_net_),
            .in3(N__24167),
            .lcout(),
            .ltout(\processor_zipi8.decode4_strobes_enables_i.un9_flag_enable_type_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_0_LC_5_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_0_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_0_LC_5_14_5 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.flag_enable_RNO_0_LC_5_14_5  (
            .in0(N__17519),
            .in1(N__23987),
            .in2(N__17513),
            .in3(N__19943),
            .lcout(),
            .ltout(\processor_zipi8.decode4_strobes_enables_i.flag_enable_type_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_LC_5_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.decode4_strobes_enables_i.flag_enable_LC_5_14_6 .LUT_INIT=16'b0000101100000000;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.flag_enable_LC_5_14_6  (
            .in0(N__21436),
            .in1(N__18928),
            .in2(N__17510),
            .in3(N__19061),
            .lcout(\processor_zipi8.flag_enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33661),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.spm_enable_LC_5_14_7 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.spm_enable_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.decode4_strobes_enables_i.spm_enable_LC_5_14_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.spm_enable_LC_5_14_7  (
            .in0(N__24168),
            .in1(N__17483),
            .in2(_gnd_net_),
            .in3(N__24315),
            .lcout(\processor_zipi8.spm_enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33661),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_0_LC_5_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_0_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.decode4alu_i.alu_mux_sel_0_LC_5_15_0 .LUT_INIT=16'b0000010000100000;
    LogicCell40 \processor_zipi8.decode4alu_i.alu_mux_sel_0_LC_5_15_0  (
            .in0(N__19870),
            .in1(N__24101),
            .in2(N__24341),
            .in3(N__21189),
            .lcout(\processor_zipi8.alu_mux_sel_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33667),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.use_zero_flag_LC_5_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.use_zero_flag_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.flags_i.use_zero_flag_LC_5_15_1 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \processor_zipi8.flags_i.use_zero_flag_LC_5_15_1  (
            .in0(N__24100),
            .in1(N__24333),
            .in2(N__21213),
            .in3(N__19871),
            .lcout(\processor_zipi8.flags_i.use_zero_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33667),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_0_LC_5_15_2 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_0_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_0_LC_5_15_2 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_0_LC_5_15_2  (
            .in0(N__33823),
            .in1(N__35745),
            .in2(N__32230),
            .in3(N__31841),
            .lcout(),
            .ltout(\processor_zipi8.alu_result_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNO_3_LC_5_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_3_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_3_LC_5_15_3 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNO_3_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__18056),
            .in2(N__18050),
            .in3(N__18043),
            .lcout(\processor_zipi8.flags_i.zero_flag_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNITLO51_LC_5_15_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNITLO51_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNITLO51_LC_5_15_4 .LUT_INIT=16'b0011110001011010;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNITLO51_LC_5_15_4  (
            .in0(N__18042),
            .in1(N__17974),
            .in2(N__19917),
            .in3(N__24099),
            .lcout(\processor_zipi8.N_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_1_LC_5_15_6 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_1_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_1_LC_5_15_6 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_1_LC_5_15_6  (
            .in0(N__33824),
            .in1(N__39127),
            .in2(N__39575),
            .in3(N__35746),
            .lcout(\processor_zipi8.alu_result_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_0_LC_5_15_7 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_0_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_0_LC_5_15_7 .LUT_INIT=16'b1100110110101011;
    LogicCell40 \processor_zipi8.decode4alu_i.arith_logical_sel_1_0_LC_5_15_7  (
            .in0(N__24098),
            .in1(N__24332),
            .in2(N__21212),
            .in3(N__19869),
            .lcout(\processor_zipi8.arith_logical_sel_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_2_LC_5_16_3 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_2_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_2_LC_5_16_3 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_2_LC_5_16_3  (
            .in0(N__33869),
            .in1(N__38310),
            .in2(N__38879),
            .in3(N__36102),
            .lcout(),
            .ltout(\processor_zipi8.alu_result_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.zero_flag_RNO_2_LC_5_16_4 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_2_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.zero_flag_RNO_2_LC_5_16_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \processor_zipi8.flags_i.zero_flag_RNO_2_LC_5_16_4  (
            .in0(N__20111),
            .in1(N__17918),
            .in2(N__17912),
            .in3(N__17909),
            .lcout(\processor_zipi8.flags_i.zero_flag_3_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__7_LC_6_1_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__7_LC_6_1_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__7_LC_6_1_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__7_LC_6_1_0  (
            .in0(N__34568),
            .in1(N__36668),
            .in2(N__33341),
            .in3(N__33015),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33680),
            .ce(N__23437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__7_LC_6_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__7_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__7_LC_6_2_0 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__7_LC_6_2_0  (
            .in0(N__34567),
            .in1(N__32980),
            .in2(N__36627),
            .in3(N__33310),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33669),
            .ce(N__22930),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__7_LC_6_3_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__7_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__7_LC_6_3_0 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__7_LC_6_3_0  (
            .in0(N__34570),
            .in1(N__32979),
            .in2(N__36803),
            .in3(N__33358),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33663),
            .ce(N__22339),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe12_0_a2_LC_6_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe12_0_a2_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe12_0_a2_LC_6_4_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe12_0_a2_LC_6_4_0  (
            .in0(N__20848),
            .in1(N__22255),
            .in2(N__23107),
            .in3(N__27392),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe20_0_a2_LC_6_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe20_0_a2_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe20_0_a2_LC_6_4_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe20_0_a2_LC_6_4_1  (
            .in0(N__27390),
            .in1(N__23099),
            .in2(N__22290),
            .in3(N__20850),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_LC_6_4_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_LC_6_4_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_LC_6_4_2  (
            .in0(N__20852),
            .in1(N__22266),
            .in2(N__23108),
            .in3(N__27394),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe4_0_a2_LC_6_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe4_0_a2_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe4_0_a2_LC_6_4_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe4_0_a2_LC_6_4_3  (
            .in0(N__27389),
            .in1(N__23103),
            .in2(N__22288),
            .in3(N__20847),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_LC_6_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_LC_6_4_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_LC_6_4_4  (
            .in0(N__20846),
            .in1(N__22251),
            .in2(N__23165),
            .in3(N__27388),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe21_0_a2_LC_6_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe21_0_a2_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe21_0_a2_LC_6_4_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe21_0_a2_LC_6_4_5  (
            .in0(N__27391),
            .in1(N__20534),
            .in2(N__22289),
            .in3(N__20849),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe6_0_a2_LC_6_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe6_0_a2_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe6_0_a2_LC_6_4_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe6_0_a2_LC_6_4_6  (
            .in0(N__23104),
            .in1(N__22262),
            .in2(N__27460),
            .in3(N__20645),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe5_0_a2_LC_6_4_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe5_0_a2_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe5_0_a2_LC_6_4_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe5_0_a2_LC_6_4_7  (
            .in0(N__27393),
            .in1(N__20535),
            .in2(N__22291),
            .in3(N__20851),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNINMK21_3_LC_6_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNINMK21_3_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNINMK21_3_LC_6_5_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNINMK21_3_LC_6_5_0  (
            .in0(N__30835),
            .in1(N__18208),
            .in2(N__31743),
            .in3(N__18194),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_bm_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI1QV11_3_LC_6_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI1QV11_3_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI1QV11_3_LC_6_5_1 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI1QV11_3_LC_6_5_1  (
            .in0(N__18161),
            .in1(N__18173),
            .in2(N__31693),
            .in3(N__30834),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_14_am_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_3_LC_6_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_3_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_3_LC_6_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_3_LC_6_5_2  (
            .in0(N__18484),
            .in1(N__18520),
            .in2(_gnd_net_),
            .in3(N__37083),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_3_LC_6_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_3_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_3_LC_6_5_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_3_LC_6_5_3  (
            .in0(N__18146),
            .in1(N__28599),
            .in2(N__18212),
            .in3(N__28924),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_3_LC_6_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_3_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_3_LC_6_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_3_LC_6_5_4  (
            .in0(N__18209),
            .in1(N__18193),
            .in2(_gnd_net_),
            .in3(N__37084),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_3_LC_6_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_3_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_3_LC_6_5_5 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_3_LC_6_5_5  (
            .in0(N__18089),
            .in1(N__18182),
            .in2(N__18176),
            .in3(N__28600),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_3_LC_6_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_3_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_3_LC_6_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_3_LC_6_5_6  (
            .in0(N__18172),
            .in1(N__18160),
            .in2(_gnd_net_),
            .in3(N__37082),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIHGK21_0_LC_6_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIHGK21_0_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIHGK21_0_LC_6_5_7 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIHGK21_0_LC_6_5_7  (
            .in0(N__18140),
            .in1(N__31718),
            .in2(N__18122),
            .in3(N__30833),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_5_LC_6_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_5_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_5_LC_6_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_5_LC_6_6_0  (
            .in0(N__37299),
            .in1(N__18307),
            .in2(_gnd_net_),
            .in3(N__18325),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_3_LC_6_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_3_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_3_LC_6_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_3_LC_6_6_1  (
            .in0(N__18349),
            .in1(N__18340),
            .in2(_gnd_net_),
            .in3(N__37298),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNILKK21_2_LC_6_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNILKK21_2_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNILKK21_2_LC_6_6_2 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNILKK21_2_LC_6_6_2  (
            .in0(N__30973),
            .in1(N__18371),
            .in2(N__18386),
            .in3(N__31581),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI0ESR1_2_LC_6_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI0ESR1_2_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI0ESR1_2_LC_6_6_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI0ESR1_2_LC_6_6_3  (
            .in0(N__31582),
            .in1(N__18461),
            .in2(N__18389),
            .in3(N__18446),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI0ESR1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_2_LC_6_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_2_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_2_LC_6_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_am_2_LC_6_6_4  (
            .in0(N__37297),
            .in1(N__18382),
            .in2(_gnd_net_),
            .in3(N__18370),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_am_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI4ISR1_3_LC_6_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI4ISR1_3_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI4ISR1_3_LC_6_6_5 .LUT_INIT=16'b1011100100110001;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI4ISR1_3_LC_6_6_5  (
            .in0(N__31583),
            .in1(N__18359),
            .in2(N__18353),
            .in3(N__18341),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI4ISR1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIRQK21_5_LC_6_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIRQK21_5_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIRQK21_5_LC_6_6_6 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIRQK21_5_LC_6_6_6  (
            .in0(N__30974),
            .in1(N__31584),
            .in2(N__18329),
            .in3(N__18308),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNICQSR1_5_LC_6_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNICQSR1_5_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNICQSR1_5_LC_6_6_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNICQSR1_5_LC_6_6_7  (
            .in0(N__31585),
            .in1(N__18295),
            .in2(N__18281),
            .in3(N__18278),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_2_LC_6_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_2_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_2_LC_6_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_am_2_LC_6_7_0  (
            .in0(N__18226),
            .in1(N__18244),
            .in2(_gnd_net_),
            .in3(N__37294),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_am_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIVNV11_2_LC_6_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIVNV11_2_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIVNV11_2_LC_6_7_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNIVNV11_2_LC_6_7_1  (
            .in0(N__18245),
            .in1(N__31390),
            .in2(N__18230),
            .in3(N__30975),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI2HMP1_2_LC_6_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI2HMP1_2_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI2HMP1_2_LC_6_7_2 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI2HMP1_2_LC_6_7_2  (
            .in0(N__31391),
            .in1(N__18557),
            .in2(N__18215),
            .in3(N__18571),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI2HMP1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_2_LC_6_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_2_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_2_LC_6_7_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_bm_2_LC_6_7_3  (
            .in0(N__37296),
            .in1(_gnd_net_),
            .in2(N__18572),
            .in3(N__18556),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_bm_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_2_LC_6_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_2_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_2_LC_6_7_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_2_LC_6_7_4  (
            .in0(N__18539),
            .in1(N__28544),
            .in2(N__18533),
            .in3(N__28955),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_2_LC_6_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_2_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_2_LC_6_7_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_2_LC_6_7_5  (
            .in0(N__28545),
            .in1(N__18425),
            .in2(N__18530),
            .in3(N__18527),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI6LMP1_3_LC_6_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI6LMP1_3_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI6LMP1_3_LC_6_7_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI6LMP1_3_LC_6_7_6  (
            .in0(N__31392),
            .in1(N__18521),
            .in2(N__18497),
            .in3(N__18485),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI6LMP1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_2_LC_6_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_2_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_2_LC_6_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_bm_2_LC_6_7_7  (
            .in0(N__37295),
            .in1(N__18457),
            .in2(_gnd_net_),
            .in3(N__18445),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIPOK21_4_LC_6_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIPOK21_4_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIPOK21_4_LC_6_8_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIPOK21_4_LC_6_8_0  (
            .in0(N__31575),
            .in1(N__18409),
            .in2(N__30942),
            .in3(N__18419),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_4_LC_6_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_4_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_4_LC_6_8_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_4_LC_6_8_1  (
            .in0(N__18418),
            .in1(N__28957),
            .in2(N__18410),
            .in3(N__37327),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_4_LC_6_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_4_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_4_LC_6_8_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_4_LC_6_8_2  (
            .in0(N__28958),
            .in1(N__18634),
            .in2(N__18392),
            .in3(N__18611),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_4_LC_6_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_4_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_4_LC_6_8_3 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_4_LC_6_8_3  (
            .in0(N__18700),
            .in1(N__18734),
            .in2(N__18686),
            .in3(N__28959),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_4_LC_6_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_4_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_4_LC_6_8_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_4_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__18743),
            .in2(N__18737),
            .in3(N__28598),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_4_LC_6_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_4_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_4_LC_6_8_5 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_4_LC_6_8_5  (
            .in0(N__18715),
            .in1(N__28956),
            .in2(N__37385),
            .in3(N__18724),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI3SV11_4_LC_6_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI3SV11_4_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI3SV11_4_LC_6_8_6 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNI3SV11_4_LC_6_8_6  (
            .in0(N__31576),
            .in1(N__31004),
            .in2(N__18728),
            .in3(N__18716),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIAPMP1_4_LC_6_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIAPMP1_4_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIAPMP1_4_LC_6_8_7 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIAPMP1_4_LC_6_8_7  (
            .in0(N__18701),
            .in1(N__18685),
            .in2(N__18665),
            .in3(N__31577),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNIAPMP1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_4_LC_6_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_4_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_4_LC_6_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_4_LC_6_9_0  (
            .in0(N__35983),
            .in1(N__18662),
            .in2(_gnd_net_),
            .in3(N__18650),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267 ),
            .ltout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__4_LC_6_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__4_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__4_LC_6_9_1 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__4_LC_6_9_1  (
            .in0(N__35340),
            .in1(N__34495),
            .in2(N__18638),
            .in3(N__35984),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33639),
            .ce(N__20287),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI8MSR1_4_LC_6_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI8MSR1_4_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI8MSR1_4_LC_6_9_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNI8MSR1_4_LC_6_9_2  (
            .in0(N__31712),
            .in1(N__18635),
            .in2(N__18620),
            .in3(N__18610),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNI8MSR1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_1_LC_6_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_1_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_1_LC_6_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_1_LC_6_9_3  (
            .in0(N__18596),
            .in1(N__18584),
            .in2(_gnd_net_),
            .in3(N__35982),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198 ),
            .ltout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__1_LC_6_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__1_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__1_LC_6_9_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram14__1_LC_6_9_4  (
            .in0(N__34494),
            .in1(N__36850),
            .in2(N__19106),
            .in3(N__39494),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33639),
            .ce(N__20287),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIS9SR1_1_LC_6_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIS9SR1_1_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIS9SR1_1_LC_6_9_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIS9SR1_1_LC_6_9_5  (
            .in0(N__20753),
            .in1(N__20732),
            .in2(N__20951),
            .in3(N__31708),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI1P541_4_LC_6_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI1P541_4_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI1P541_4_LC_6_9_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI1P541_4_LC_6_9_6  (
            .in0(N__30917),
            .in1(N__24953),
            .in2(N__31741),
            .in3(N__25109),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_4_LC_6_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_4_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_4_LC_6_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_4_LC_6_9_7  (
            .in0(N__24952),
            .in1(N__25108),
            .in2(_gnd_net_),
            .in3(N__37429),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_3_LC_6_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_3_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_3_LC_6_10_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_3_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__19103),
            .in2(_gnd_net_),
            .in3(N__19085),
            .lcout(\processor_zipi8.arith_logical_result_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33646),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_0_LC_6_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_0_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_0_LC_6_10_1 .LUT_INIT=16'b0000111000001010;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.register_enable_RNO_0_LC_6_10_1  (
            .in0(N__18925),
            .in1(N__19963),
            .in2(N__19079),
            .in3(N__24166),
            .lcout(),
            .ltout(\processor_zipi8.decode4_strobes_enables_i.register_enable_type_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_LC_6_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.decode4_strobes_enables_i.register_enable_LC_6_10_2 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.register_enable_LC_6_10_2  (
            .in0(N__21391),
            .in1(N__19031),
            .in2(N__18935),
            .in3(N__18926),
            .lcout(\processor_zipi8.register_enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33646),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_4_LC_6_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_4_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_4_LC_6_10_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_4_LC_6_10_3  (
            .in0(N__18812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19258),
            .lcout(\processor_zipi8.arith_logical_result_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33646),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical4_process_carry_arith_logical_28_4_LC_6_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical4_process_carry_arith_logical_28_4_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical4_process_carry_arith_logical_28_4_LC_6_10_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical4_process_carry_arith_logical_28_4_LC_6_10_4  (
            .in0(N__19776),
            .in1(N__21846),
            .in2(N__19259),
            .in3(N__18811),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4 ),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_28_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical5_process_carry_arith_logical_34_5_LC_6_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical5_process_carry_arith_logical_34_5_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical5_process_carry_arith_logical_34_5_LC_6_10_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.calc_carry_arith_logical5_process_carry_arith_logical_34_5_LC_6_10_5  (
            .in0(N__18797),
            .in1(N__19321),
            .in2(N__19334),
            .in3(N__19777),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.carry_arith_logical_34_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_5_LC_6_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_5_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_5_LC_6_10_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.arith_logical_result_5_LC_6_10_6  (
            .in0(N__19322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19310),
            .lcout(\processor_zipi8.arith_logical_result_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33646),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.flags_i.carry_flag_RNO_6_LC_6_10_7 .C_ON=1'b0;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_6_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.flags_i.carry_flag_RNO_6_LC_6_10_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \processor_zipi8.flags_i.carry_flag_RNO_6_LC_6_10_7  (
            .in0(N__35297),
            .in1(N__37899),
            .in2(N__38731),
            .in3(N__30207),
            .lcout(\processor_zipi8.flags_i.parity_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_LC_6_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_LC_6_11_0 .LUT_INIT=16'b1011101100000101;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_LC_6_11_0  (
            .in0(N__21683),
            .in1(N__23989),
            .in2(N__19556),
            .in3(N__19499),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_LC_6_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_LC_6_11_1 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_LC_6_11_1  (
            .in0(N__19397),
            .in1(N__21684),
            .in2(N__19298),
            .in3(N__19295),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tz_4_LC_6_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tz_4_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tz_4_LC_6_11_2 .LUT_INIT=16'b0000111110111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tz_4_LC_6_11_2  (
            .in0(N__19203),
            .in1(N__21821),
            .in2(N__19782),
            .in3(N__19472),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_tzZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_4_LC_6_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_4_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_4_LC_6_11_3 .LUT_INIT=16'b0011111000000010;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_4_LC_6_11_3  (
            .in0(N__23990),
            .in1(N__19234),
            .in2(N__21836),
            .in3(N__19536),
            .lcout(),
            .ltout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_LC_6_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_LC_6_11_4 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_4_LC_6_11_4  (
            .in0(N__19236),
            .in1(N__19268),
            .in2(N__19262),
            .in3(N__19112),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_4_LC_6_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_4_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_4_LC_6_11_5 .LUT_INIT=16'b0100001101111111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1_4_LC_6_11_5  (
            .in0(N__19471),
            .in1(N__19235),
            .in2(N__21835),
            .in3(N__19204),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_1_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_1_LC_6_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_1_LC_6_11_6 .LUT_INIT=16'b0010001001011111;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1_1_LC_6_11_6  (
            .in0(N__21682),
            .in1(N__19617),
            .in2(N__19555),
            .in3(N__21546),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_3_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_1_LC_6_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_1_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_1_LC_6_11_7 .LUT_INIT=16'b0101110111011101;
    LogicCell40 \processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_1_LC_6_11_7  (
            .in0(N__21547),
            .in1(N__19493),
            .in2(N__19482),
            .in3(N__19751),
            .lcout(\processor_zipi8.arith_and_logic_operations_i.half_arith_logical_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNINIG61_4_LC_6_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNINIG61_4_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNINIG61_4_LC_6_12_0 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNINIG61_4_LC_6_12_0  (
            .in0(N__31009),
            .in1(N__19376),
            .in2(N__32528),
            .in3(N__31573),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI4AK32_4_LC_6_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI4AK32_4_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI4AK32_4_LC_6_12_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI4AK32_4_LC_6_12_1  (
            .in0(N__31574),
            .in1(N__23359),
            .in2(N__19391),
            .in3(N__33731),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI4AK32_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_4_LC_6_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_4_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_4_LC_6_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_4_LC_6_12_2  (
            .in0(N__37424),
            .in1(N__22978),
            .in2(_gnd_net_),
            .in3(N__27707),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_4_LC_6_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_4_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_4_LC_6_12_3 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_4_LC_6_12_3  (
            .in0(N__28647),
            .in1(N__19388),
            .in2(N__19379),
            .in3(N__29001),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_4_LC_6_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_4_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_4_LC_6_12_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_4_LC_6_12_4  (
            .in0(N__37425),
            .in1(_gnd_net_),
            .in2(N__23360),
            .in3(N__33730),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_4_LC_6_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_4_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_4_LC_6_12_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_4_LC_6_12_5  (
            .in0(N__19375),
            .in1(N__32524),
            .in2(_gnd_net_),
            .in3(N__37426),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_4_LC_6_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_4_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_4_LC_6_12_6 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_4_LC_6_12_6  (
            .in0(N__19358),
            .in1(N__19352),
            .in2(N__19346),
            .in3(N__28648),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_4_LC_6_12_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_4_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_4_LC_6_12_7 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_4_LC_6_12_7  (
            .in0(N__25603),
            .in1(N__19979),
            .in2(N__25160),
            .in3(N__25763),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_2_LC_6_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_2_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4alu_i.arith_logical_sel_1_2_LC_6_13_0 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \processor_zipi8.decode4alu_i.arith_logical_sel_1_2_LC_6_13_0  (
            .in0(N__19918),
            .in1(N__24310),
            .in2(_gnd_net_),
            .in3(N__24126),
            .lcout(\processor_zipi8.arith_logical_sel_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_3_LC_6_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_3_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_3_LC_6_13_2 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_3_LC_6_13_2  (
            .in0(N__28646),
            .in1(N__23579),
            .in2(N__20153),
            .in3(N__19664),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_3_LC_6_13_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_3_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_3_LC_6_13_3 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_3_LC_6_13_3  (
            .in0(N__25601),
            .in1(N__19682),
            .in2(N__19670),
            .in3(N__25762),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_3_LC_6_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_3_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_3_LC_6_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_3_LC_6_13_4  (
            .in0(N__21931),
            .in1(N__23485),
            .in2(_gnd_net_),
            .in3(N__37423),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_3_LC_6_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_3_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_3_LC_6_13_5 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_3_LC_6_13_5  (
            .in0(N__25970),
            .in1(N__28645),
            .in2(N__19667),
            .in3(N__28997),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_3_LC_6_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_3_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_3_LC_6_13_6 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_3_LC_6_13_6  (
            .in0(N__27821),
            .in1(N__25602),
            .in2(N__26267),
            .in3(N__19658),
            .lcout(\processor_zipi8.sy_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIPPE01_3_LC_6_14_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIPPE01_3_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIPPE01_3_LC_6_14_0 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIPPE01_3_LC_6_14_0  (
            .in0(N__31008),
            .in1(N__23600),
            .in2(N__23621),
            .in3(N__31572),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_bm_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI8OGN1_3_LC_6_14_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI8OGN1_3_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI8OGN1_3_LC_6_14_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI8OGN1_3_LC_6_14_1  (
            .in0(N__20165),
            .in1(N__22388),
            .in2(N__19643),
            .in3(N__31570),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI8OGN1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU6AG4_3_LC_6_14_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU6AG4_3_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU6AG4_3_LC_6_14_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIU6AG4_3_LC_6_14_2  (
            .in0(N__20099),
            .in1(N__27312),
            .in2(N__20105),
            .in3(N__27609),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIHPTE1_3_LC_6_14_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIHPTE1_3_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIHPTE1_3_LC_6_14_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIHPTE1_3_LC_6_14_3  (
            .in0(N__21932),
            .in1(N__31569),
            .in2(N__23486),
            .in3(N__31007),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_7_am_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIONE42_3_LC_6_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIONE42_3_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIONE42_3_LC_6_14_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIONE42_3_LC_6_14_4  (
            .in0(N__26207),
            .in1(N__25985),
            .in2(N__20102),
            .in3(N__31571),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIONE42_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINP2G8_3_LC_6_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINP2G8_3_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINP2G8_3_LC_6_14_5 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINP2G8_3_LC_6_14_5  (
            .in0(N__27313),
            .in1(N__20093),
            .in2(N__20081),
            .in3(N__20066),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNINP2G8_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5OSHH_3_LC_6_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5OSHH_3_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5OSHH_3_LC_6_14_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5OSHH_3_LC_6_14_6  (
            .in0(N__22169),
            .in1(N__27110),
            .in2(N__20060),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.sx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__0_LC_6_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__0_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__0_LC_6_15_0 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__0_LC_6_15_0  (
            .in0(N__35976),
            .in1(N__33903),
            .in2(N__32289),
            .in3(N__31997),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33679),
            .ce(N__20140),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__1_LC_6_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__1_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__1_LC_6_15_1 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__1_LC_6_15_1  (
            .in0(N__33902),
            .in1(N__39544),
            .in2(N__39227),
            .in3(N__35981),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33679),
            .ce(N__20140),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__2_LC_6_15_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__2_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__2_LC_6_15_2 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__2_LC_6_15_2  (
            .in0(N__35977),
            .in1(N__38847),
            .in2(N__34276),
            .in3(N__38446),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33679),
            .ce(N__20140),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_2_LC_6_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_2_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_2_LC_6_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_2_LC_6_15_3  (
            .in0(N__22399),
            .in1(N__21790),
            .in2(_gnd_net_),
            .in3(N__37503),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__3_LC_6_15_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__3_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__3_LC_6_15_4 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__3_LC_6_15_4  (
            .in0(N__35978),
            .in1(N__33904),
            .in2(N__38159),
            .in3(N__37627),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33679),
            .ce(N__20140),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_3_LC_6_15_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_3_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_3_LC_6_15_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_3_LC_6_15_5  (
            .in0(N__22387),
            .in1(N__20164),
            .in2(_gnd_net_),
            .in3(N__37504),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__4_LC_6_15_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__4_LC_6_15_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__4_LC_6_15_6 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__4_LC_6_15_6  (
            .in0(N__35979),
            .in1(N__35347),
            .in2(N__35097),
            .in3(N__33908),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33679),
            .ce(N__20140),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__5_LC_6_15_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__5_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__5_LC_6_15_7 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__5_LC_6_15_7  (
            .in0(N__30089),
            .in1(N__35980),
            .in2(N__34078),
            .in3(N__30390),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33679),
            .ce(N__20140),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_4_LC_6_16_2 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_4_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_4_LC_6_16_2 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_3_4_LC_6_16_2  (
            .in0(N__33825),
            .in1(N__35007),
            .in2(N__35413),
            .in3(N__36101),
            .lcout(\processor_zipi8.alu_result_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__7_LC_7_1_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__7_LC_7_1_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__7_LC_7_1_0 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__7_LC_7_1_0  (
            .in0(N__34325),
            .in1(N__33002),
            .in2(N__36792),
            .in3(N__33327),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33690),
            .ce(N__27781),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__5_LC_7_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__5_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__5_LC_7_2_0 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__5_LC_7_2_0  (
            .in0(N__30464),
            .in1(N__34580),
            .in2(N__30134),
            .in3(N__36625),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33682),
            .ce(N__32497),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__6_LC_7_2_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__6_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__6_LC_7_2_1 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__6_LC_7_2_1  (
            .in0(N__34579),
            .in1(N__36623),
            .in2(N__29782),
            .in3(N__29291),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33682),
            .ce(N__32497),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__7_LC_7_2_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__7_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__7_LC_7_2_2 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__7_LC_7_2_2  (
            .in0(N__33301),
            .in1(N__36624),
            .in2(N__33010),
            .in3(N__34581),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33682),
            .ce(N__32497),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI7V541_7_LC_7_3_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI7V541_7_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI7V541_7_LC_7_3_0 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI7V541_7_LC_7_3_0  (
            .in0(N__20186),
            .in1(N__31734),
            .in2(N__31022),
            .in3(N__21581),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI43VU1_7_LC_7_3_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI43VU1_7_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI43VU1_7_LC_7_3_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI43VU1_7_LC_7_3_1  (
            .in0(N__31735),
            .in1(N__20203),
            .in2(N__20237),
            .in3(N__22577),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI43VU1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNITOG61_7_LC_7_3_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNITOG61_7_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNITOG61_7_LC_7_3_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNITOG61_7_LC_7_3_2  (
            .in0(N__21607),
            .in1(N__31736),
            .in2(N__32714),
            .in3(N__31013),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIGMK32_7_LC_7_3_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIGMK32_7_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIGMK32_7_LC_7_3_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIGMK32_7_LC_7_3_3  (
            .in0(N__31737),
            .in1(N__23315),
            .in2(N__20234),
            .in3(N__23872),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIGMK32_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIGUM4_7_LC_7_3_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIGUM4_7_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIGUM4_7_LC_7_3_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIGUM4_7_LC_7_3_4  (
            .in0(N__20231),
            .in1(N__27286),
            .in2(N__20225),
            .in3(N__27629),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_7_LC_7_3_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_7_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_7_LC_7_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_7_LC_7_3_5  (
            .in0(N__20204),
            .in1(N__22576),
            .in2(_gnd_net_),
            .in3(N__37355),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_7_LC_7_3_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_7_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_7_LC_7_3_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_7_LC_7_3_6  (
            .in0(N__20171),
            .in1(N__28658),
            .in2(N__20189),
            .in3(N__28968),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_7_LC_7_3_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_7_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_7_LC_7_3_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_7_LC_7_3_7  (
            .in0(N__21580),
            .in1(N__20185),
            .in2(_gnd_net_),
            .in3(N__37354),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe31_0_a2_LC_7_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe31_0_a2_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe31_0_a2_LC_7_4_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe31_0_a2_LC_7_4_0  (
            .in0(N__20642),
            .in1(N__22268),
            .in2(N__20541),
            .in3(N__27430),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe19_0_a2_LC_7_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe19_0_a2_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe19_0_a2_LC_7_4_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe19_0_a2_LC_7_4_1  (
            .in0(N__27428),
            .in1(N__20332),
            .in2(N__22292),
            .in3(N__20639),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe7_0_a2_LC_7_4_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe7_0_a2_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe7_0_a2_LC_7_4_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe7_0_a2_LC_7_4_2  (
            .in0(N__20644),
            .in1(N__22267),
            .in2(N__20542),
            .in3(N__27429),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe3_0_a2_LC_7_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe3_0_a2_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe3_0_a2_LC_7_4_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe3_0_a2_LC_7_4_3  (
            .in0(N__27433),
            .in1(N__20333),
            .in2(N__22294),
            .in3(N__20643),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe14_0_a2_LC_7_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe14_0_a2_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe14_0_a2_LC_7_4_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe14_0_a2_LC_7_4_4  (
            .in0(N__20638),
            .in1(N__22279),
            .in2(N__23105),
            .in3(N__27435),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe22_0_a2_LC_7_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe22_0_a2_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe22_0_a2_LC_7_4_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe22_0_a2_LC_7_4_5  (
            .in0(N__27432),
            .in1(N__23092),
            .in2(N__22293),
            .in3(N__20640),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe30_0_a2_LC_7_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe30_0_a2_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe30_0_a2_LC_7_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe30_0_a2_LC_7_4_6  (
            .in0(N__20641),
            .in1(N__22272),
            .in2(N__23106),
            .in3(N__27431),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_LC_7_4_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_LC_7_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_LC_7_4_7  (
            .in0(N__27434),
            .in1(N__20527),
            .in2(N__22295),
            .in3(N__20853),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI7JI91_4_LC_7_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI7JI91_4_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI7JI91_4_LC_7_5_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI7JI91_4_LC_7_5_0  (
            .in0(N__30822),
            .in1(N__26075),
            .in2(N__31703),
            .in3(N__24521),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNII4IQ1_4_LC_7_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNII4IQ1_4_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNII4IQ1_4_LC_7_5_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNII4IQ1_4_LC_7_5_1  (
            .in0(N__24482),
            .in1(N__24499),
            .in2(N__20258),
            .in3(N__31623),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNII4IQ1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNI12F01_7_LC_7_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNI12F01_7_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNI12F01_7_LC_7_5_2 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNI12F01_7_LC_7_5_2  (
            .in0(N__30823),
            .in1(N__20489),
            .in2(N__31704),
            .in3(N__20468),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIO8HN1_7_LC_7_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIO8HN1_7_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIO8HN1_7_LC_7_5_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIO8HN1_7_LC_7_5_3  (
            .in0(N__20440),
            .in1(N__20426),
            .in2(N__20255),
            .in3(N__31624),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNIO8HN1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_7_LC_7_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_7_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_7_LC_7_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_7_LC_7_5_4  (
            .in0(N__20485),
            .in1(N__20467),
            .in2(_gnd_net_),
            .in3(N__37214),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_7_LC_7_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_7_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_7_LC_7_5_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_7_LC_7_5_5  (
            .in0(N__37215),
            .in1(_gnd_net_),
            .in2(N__20441),
            .in3(N__20425),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIJJE01_0_LC_7_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIJJE01_0_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIJJE01_0_LC_7_5_6 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIJJE01_0_LC_7_5_6  (
            .in0(N__31616),
            .in1(N__23276),
            .in2(N__30921),
            .in3(N__23411),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe24_0_a2_LC_7_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe24_0_a2_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe24_0_a2_LC_7_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe24_0_a2_LC_7_5_7  (
            .in0(N__20831),
            .in1(N__27289),
            .in2(N__22283),
            .in3(N__23146),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.awe24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_5_LC_7_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_5_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_5_LC_7_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_5_LC_7_6_0  (
            .in0(N__37332),
            .in1(N__29812),
            .in2(_gnd_net_),
            .in3(N__22648),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_5_LC_7_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_5_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_5_LC_7_6_1 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_5_LC_7_6_1  (
            .in0(N__20339),
            .in1(N__20666),
            .in2(N__20402),
            .in3(N__28602),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIO5SR1_0_LC_7_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIO5SR1_0_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIO5SR1_0_LC_7_6_2 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram15__RNIO5SR1_0_LC_7_6_2  (
            .in0(N__20386),
            .in1(N__20369),
            .in2(N__20348),
            .in3(N__31713),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram15__RNIO5SR1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_5_LC_7_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_5_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_5_LC_7_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_5_LC_7_6_3  (
            .in0(N__22948),
            .in1(N__22747),
            .in2(_gnd_net_),
            .in3(N__37328),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_5_LC_7_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_5_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_5_LC_7_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_5_LC_7_6_4  (
            .in0(N__37330),
            .in1(N__23338),
            .in2(_gnd_net_),
            .in3(N__23890),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_5_LC_7_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_5_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_5_LC_7_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_5_LC_7_6_5  (
            .in0(N__22768),
            .in1(N__24940),
            .in2(_gnd_net_),
            .in3(N__37329),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_5_LC_7_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_5_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_5_LC_7_6_6 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_5_LC_7_6_6  (
            .in0(N__28601),
            .in1(N__20675),
            .in2(N__20669),
            .in3(N__28885),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_6_LC_7_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_6_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_6_LC_7_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_6_LC_7_6_7  (
            .in0(N__29095),
            .in1(N__22442),
            .in2(_gnd_net_),
            .in3(N__37331),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_2_LC_7_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_2_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_2_LC_7_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_2_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__20873),
            .in2(_gnd_net_),
            .in3(N__31428),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIBJTE1_0_LC_7_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIBJTE1_0_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIBJTE1_0_LC_7_7_1 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIBJTE1_0_LC_7_7_1  (
            .in0(N__31425),
            .in1(N__23534),
            .in2(N__31017),
            .in3(N__21979),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNICBE42_0_LC_7_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNICBE42_0_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNICBE42_0_LC_7_7_2 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNICBE42_0_LC_7_7_2  (
            .in0(N__25448),
            .in1(N__25913),
            .in2(N__20582),
            .in3(N__31426),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNICBE42_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6E9G4_0_LC_7_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6E9G4_0_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6E9G4_0_LC_7_7_3 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6E9G4_0_LC_7_7_3  (
            .in0(N__27287),
            .in1(N__27594),
            .in2(N__20579),
            .in3(N__20768),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI781G8_0_LC_7_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI781G8_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI781G8_0_LC_7_7_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI781G8_0_LC_7_7_4  (
            .in0(N__27288),
            .in1(N__20576),
            .in2(N__20564),
            .in3(N__20561),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI781G8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_0_LC_7_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_0_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_0_LC_7_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe29_0_a2_0_LC_7_7_5  (
            .in0(N__31000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27595),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_1_LC_7_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_1_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_1_LC_7_7_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe0_0_a2_1_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__20872),
            .in2(_gnd_net_),
            .in3(N__31427),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNISBGN1_0_LC_7_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNISBGN1_0_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNISBGN1_0_LC_7_7_7 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNISBGN1_0_LC_7_7_7  (
            .in0(N__31424),
            .in1(N__20900),
            .in2(N__21920),
            .in3(N__20777),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNISBGN1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIUCMP1_1_LC_7_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIUCMP1_1_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIUCMP1_1_LC_7_8_0 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNIUCMP1_1_LC_7_8_0  (
            .in0(N__31707),
            .in1(N__21017),
            .in2(N__20762),
            .in3(N__20999),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNITLV11_1_LC_7_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNITLV11_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNITLV11_1_LC_7_8_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram9__RNITLV11_1_LC_7_8_1  (
            .in0(N__20714),
            .in1(N__31706),
            .in2(N__20696),
            .in3(N__30848),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_10_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_1_LC_7_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_1_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_1_LC_7_8_2 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_1_LC_7_8_2  (
            .in0(N__37323),
            .in1(N__20965),
            .in2(N__28998),
            .in3(N__20980),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_LC_7_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_LC_7_8_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_13_ns_1_LC_7_8_3  (
            .in0(N__20752),
            .in1(N__20731),
            .in2(N__20720),
            .in3(N__28954),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_13_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_LC_7_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_LC_7_8_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_14_ns_1_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__20987),
            .in2(N__20717),
            .in3(N__28587),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_14_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_1_LC_7_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_1_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_1_LC_7_8_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_1_LC_7_8_5  (
            .in0(N__20713),
            .in1(N__28949),
            .in2(N__20695),
            .in3(N__37322),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_LC_7_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_LC_7_8_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_10_ns_1_LC_7_8_6  (
            .in0(N__28950),
            .in1(N__21016),
            .in2(N__21002),
            .in3(N__20998),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_10_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIJIK21_1_LC_7_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIJIK21_1_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIJIK21_1_LC_7_8_7 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram12__RNIJIK21_1_LC_7_8_7  (
            .in0(N__20981),
            .in1(N__31705),
            .in2(N__20969),
            .in3(N__30847),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_13_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_7_LC_7_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_7_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_7_LC_7_9_0 .LUT_INIT=16'b1101100001010101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_7_LC_7_9_0  (
            .in0(N__20942),
            .in1(N__21587),
            .in2(N__20912),
            .in3(N__28586),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_0_LC_7_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_0_LC_7_9_1 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_0_LC_7_9_1  (
            .in0(N__28927),
            .in1(N__37301),
            .in2(N__21980),
            .in3(N__23533),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_0_LC_7_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_0_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_0_LC_7_9_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_0_LC_7_9_2  (
            .in0(N__28929),
            .in1(N__25912),
            .in2(N__20918),
            .in3(N__25447),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_0_LC_7_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_0_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_0_LC_7_9_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_0_LC_7_9_3  (
            .in0(N__28585),
            .in1(_gnd_net_),
            .in2(N__20915),
            .in3(N__20879),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_7_LC_7_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_7_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_7_LC_7_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_7_LC_7_9_4  (
            .in0(N__37303),
            .in1(N__23311),
            .in2(_gnd_net_),
            .in3(N__23873),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_0_LC_7_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_0_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_0_LC_7_9_5 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_0_LC_7_9_5  (
            .in0(N__28926),
            .in1(N__37300),
            .in2(N__23275),
            .in3(N__23407),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_0_LC_7_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_0_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_0_LC_7_9_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_0_LC_7_9_6  (
            .in0(N__28928),
            .in1(N__21913),
            .in2(N__20903),
            .in3(N__20896),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_7_LC_7_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_7_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_7_LC_7_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_7_LC_7_9_7  (
            .in0(N__32701),
            .in1(N__21608),
            .in2(_gnd_net_),
            .in3(N__37302),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__5_LC_7_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__5_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__5_LC_7_10_0 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__5_LC_7_10_0  (
            .in0(N__30034),
            .in1(N__36525),
            .in2(N__34824),
            .in3(N__30269),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33650),
            .ce(N__25091),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__6_LC_7_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__6_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__6_LC_7_10_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__6_LC_7_10_1  (
            .in0(N__36524),
            .in1(N__29642),
            .in2(N__29397),
            .in3(N__34711),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33650),
            .ce(N__25091),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__7_LC_7_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__7_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__7_LC_7_10_2 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__7_LC_7_10_2  (
            .in0(N__32823),
            .in1(N__36526),
            .in2(N__34825),
            .in3(N__33219),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33650),
            .ce(N__25091),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_6_0_LC_7_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_6_0_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_6_0_LC_7_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.sel_of_2nd_op_to_alu_and_port_id_i.un1_sy_6_0_LC_7_10_3  (
            .in0(N__21507),
            .in1(N__21389),
            .in2(_gnd_net_),
            .in3(N__23191),
            .lcout(\processor_zipi8.port_id_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI7UF21_1_LC_7_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI7UF21_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI7UF21_1_LC_7_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNI7UF21_1_LC_7_10_4  (
            .in0(N__21388),
            .in1(N__21533),
            .in2(_gnd_net_),
            .in3(N__21508),
            .lcout(\processor_zipi8.pc_vector_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIC1G21_4_LC_7_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIC1G21_4_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIC1G21_4_LC_7_10_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_RNIC1G21_4_LC_7_10_5  (
            .in0(N__21470),
            .in1(N__21390),
            .in2(_gnd_net_),
            .in3(N__37427),
            .lcout(\processor_zipi8.pc_vector_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.sel_of_out_port_value_i.un1_sx_7_0_LC_7_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.sel_of_out_port_value_i.un1_sx_7_0_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.sel_of_out_port_value_i.un1_sx_7_0_LC_7_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.sel_of_out_port_value_i.un1_sx_7_0_LC_7_10_6  (
            .in0(N__37428),
            .in1(N__21226),
            .in2(_gnd_net_),
            .in3(N__21110),
            .lcout(LED1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNILLE01_1_LC_7_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNILLE01_1_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNILLE01_1_LC_7_11_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNILLE01_1_LC_7_11_0  (
            .in0(N__30945),
            .in1(N__25405),
            .in2(N__31568),
            .in3(N__25424),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI0GGN1_1_LC_7_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI0GGN1_1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI0GGN1_1_LC_7_11_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI0GGN1_1_LC_7_11_1  (
            .in0(N__25370),
            .in1(N__25391),
            .in2(N__21755),
            .in3(N__31398),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_119_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIEM9G4_1_LC_7_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIEM9G4_1_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIEM9G4_1_LC_7_11_2 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIEM9G4_1_LC_7_11_2  (
            .in0(N__27277),
            .in1(N__21746),
            .in2(N__21752),
            .in3(N__27564),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIDLTE1_1_LC_7_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIDLTE1_1_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIDLTE1_1_LC_7_11_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIDLTE1_1_LC_7_11_3  (
            .in0(N__23249),
            .in1(N__31393),
            .in2(N__23510),
            .in3(N__30944),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIGFE42_1_LC_7_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIGFE42_1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIGFE42_1_LC_7_11_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIGFE42_1_LC_7_11_4  (
            .in0(N__31394),
            .in1(N__25883),
            .in2(N__21749),
            .in3(N__26033),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINO1G8_1_LC_7_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINO1G8_1_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINO1G8_1_LC_7_11_5 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNINO1G8_1_LC_7_11_5  (
            .in0(N__21740),
            .in1(N__27278),
            .in2(N__21731),
            .in3(N__21716),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_191_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5MQHH_1_LC_7_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5MQHH_1_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5MQHH_1_LC_7_11_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5MQHH_1_LC_7_11_6  (
            .in0(N__22159),
            .in1(_gnd_net_),
            .in2(N__21710),
            .in3(N__26477),
            .lcout(\processor_zipi8.sx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFIBI8_4_LC_7_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFIBI8_4_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFIBI8_4_LC_7_12_0 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFIBI8_4_LC_7_12_0  (
            .in0(N__26666),
            .in1(N__21614),
            .in2(N__21650),
            .in3(N__27275),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFIBI8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIOMUU1_4_LC_7_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIOMUU1_4_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIOMUU1_4_LC_7_12_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIOMUU1_4_LC_7_12_1  (
            .in0(N__22979),
            .in1(N__27706),
            .in2(N__21638),
            .in3(N__31688),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIOMUU1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQNTM4_4_LC_7_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQNTM4_4_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQNTM4_4_LC_7_12_2 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQNTM4_4_LC_7_12_2  (
            .in0(N__21623),
            .in1(N__27273),
            .in2(N__21617),
            .in3(N__27610),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7A3G8_4_LC_7_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7A3G8_4_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7A3G8_4_LC_7_12_3 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI7A3G8_4_LC_7_12_3  (
            .in0(N__27276),
            .in1(N__21896),
            .in2(N__21884),
            .in3(N__21803),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI7A3G8_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5PTHH_4_LC_7_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5PTHH_4_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5PTHH_4_LC_7_12_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5PTHH_4_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__21869),
            .in2(N__21863),
            .in3(N__22231),
            .lcout(\processor_zipi8.sx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNISRE42_4_LC_7_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNISRE42_4_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNISRE42_4_LC_7_12_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNISRE42_4_LC_7_12_5  (
            .in0(N__26189),
            .in1(N__25283),
            .in2(N__25121),
            .in3(N__31689),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNISRE42_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6FAG4_4_LC_7_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6FAG4_4_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6FAG4_4_LC_7_12_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI6FAG4_4_LC_7_12_6  (
            .in0(N__23177),
            .in1(N__27274),
            .in2(N__21806),
            .in3(N__27611),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIFNTE1_2_LC_7_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIFNTE1_2_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIFNTE1_2_LC_7_13_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIFNTE1_2_LC_7_13_0  (
            .in0(N__25489),
            .in1(N__31512),
            .in2(N__25508),
            .in3(N__31006),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNINNE01_2_LC_7_13_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNINNE01_2_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNINNE01_2_LC_7_13_1 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNINNE01_2_LC_7_13_1  (
            .in0(N__31005),
            .in1(N__23387),
            .in2(N__31673),
            .in3(N__23375),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI4KGN1_2_LC_7_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI4KGN1_2_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI4KGN1_2_LC_7_13_2 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNI4KGN1_2_LC_7_13_2  (
            .in0(N__22403),
            .in1(N__21797),
            .in2(N__21779),
            .in3(N__31513),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNI4KGN1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIKJE42_2_LC_7_13_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIKJE42_2_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIKJE42_2_LC_7_13_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIKJE42_2_LC_7_13_3  (
            .in0(N__31514),
            .in1(N__25859),
            .in2(N__21776),
            .in3(N__26009),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram2__RNIKJE42_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMU9G4_2_LC_7_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMU9G4_2_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMU9G4_2_LC_7_13_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIMU9G4_2_LC_7_13_4  (
            .in0(N__21767),
            .in1(N__27314),
            .in2(N__21758),
            .in3(N__27605),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI792G8_2_LC_7_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI792G8_2_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI792G8_2_LC_7_13_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram11__RNI792G8_2_LC_7_13_5  (
            .in0(N__27315),
            .in1(N__22328),
            .in2(N__22313),
            .in3(N__22310),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram11__RNI792G8_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5NRHH_2_LC_7_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5NRHH_2_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5NRHH_2_LC_7_13_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI5NRHH_2_LC_7_13_6  (
            .in0(N__22230),
            .in1(_gnd_net_),
            .in2(N__22052),
            .in3(N__27041),
            .lcout(\processor_zipi8.sx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__0_LC_7_14_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__0_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__0_LC_7_14_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__0_LC_7_14_0  (
            .in0(N__34826),
            .in1(N__32264),
            .in2(N__32027),
            .in3(N__35847),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33681),
            .ce(N__25346),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__2_LC_7_14_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__2_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__2_LC_7_14_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__2_LC_7_14_3  (
            .in0(N__35844),
            .in1(N__38830),
            .in2(N__38506),
            .in3(N__34828),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33681),
            .ce(N__25346),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_3_LC_7_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_3_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_3_LC_7_14_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_3_LC_7_14_4  (
            .in0(N__21962),
            .in1(N__21950),
            .in2(_gnd_net_),
            .in3(N__35843),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266 ),
            .ltout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__3_LC_7_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__3_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__3_LC_7_14_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__3_LC_7_14_5  (
            .in0(N__35845),
            .in1(N__38071),
            .in2(N__21935),
            .in3(N__34830),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33681),
            .ce(N__25346),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__1_LC_7_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__1_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__1_LC_7_14_6 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__1_LC_7_14_6  (
            .in0(N__34827),
            .in1(N__39178),
            .in2(N__39635),
            .in3(N__35848),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33681),
            .ce(N__25346),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__5_LC_7_14_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__5_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__5_LC_7_14_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__5_LC_7_14_7  (
            .in0(N__35846),
            .in1(N__34829),
            .in2(N__30490),
            .in3(N__30024),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33681),
            .ce(N__25346),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__0_LC_7_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__0_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__0_LC_7_15_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__0_LC_7_15_0  (
            .in0(N__34068),
            .in1(N__35973),
            .in2(N__32403),
            .in3(N__32022),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33689),
            .ce(N__22352),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__1_LC_7_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__1_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__1_LC_7_15_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__1_LC_7_15_1  (
            .in0(N__35969),
            .in1(N__34071),
            .in2(N__39644),
            .in3(N__39225),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33689),
            .ce(N__22352),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__2_LC_7_15_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__2_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__2_LC_7_15_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__2_LC_7_15_2  (
            .in0(N__34069),
            .in1(N__35975),
            .in2(N__38518),
            .in3(N__38874),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33689),
            .ce(N__22352),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__3_LC_7_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__3_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__3_LC_7_15_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__3_LC_7_15_3  (
            .in0(N__35970),
            .in1(N__38144),
            .in2(N__37706),
            .in3(N__34073),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33689),
            .ce(N__22352),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__4_LC_7_15_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__4_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__4_LC_7_15_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__4_LC_7_15_4  (
            .in0(N__34070),
            .in1(N__35974),
            .in2(N__35230),
            .in3(N__35530),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33689),
            .ce(N__22352),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__5_LC_7_15_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__5_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__5_LC_7_15_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__5_LC_7_15_5  (
            .in0(N__35971),
            .in1(N__30485),
            .in2(N__30088),
            .in3(N__34074),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33689),
            .ce(N__22352),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_5_LC_7_15_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_5_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_5_LC_7_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_bm_5_LC_7_15_6  (
            .in0(N__23704),
            .in1(N__23686),
            .in2(_gnd_net_),
            .in3(N__37487),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__6_LC_7_15_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__6_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__6_LC_7_15_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram7__6_LC_7_15_7  (
            .in0(N__35972),
            .in1(N__34072),
            .in2(N__29773),
            .in3(N__29396),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33689),
            .ce(N__22352),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__6_LC_8_1_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__6_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__6_LC_8_1_0 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__6_LC_8_1_0  (
            .in0(N__34326),
            .in1(N__29447),
            .in2(N__36793),
            .in3(N__29735),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33701),
            .ce(N__24413),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__5_LC_8_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__5_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__5_LC_8_2_0 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__5_LC_8_2_0  (
            .in0(N__34796),
            .in1(N__36656),
            .in2(N__30146),
            .in3(N__30500),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33692),
            .ce(N__27679),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__6_LC_8_2_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__6_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__6_LC_8_2_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__6_LC_8_2_1  (
            .in0(N__36655),
            .in1(N__34798),
            .in2(N__29783),
            .in3(N__29445),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33692),
            .ce(N__27679),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__7_LC_8_2_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__7_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__7_LC_8_2_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__7_LC_8_2_2  (
            .in0(N__34797),
            .in1(N__36657),
            .in2(N__33021),
            .in3(N__33302),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33692),
            .ce(N__27679),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_6_LC_8_2_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_6_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_6_LC_8_2_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_6_LC_8_2_3  (
            .in0(N__22592),
            .in1(N__22609),
            .in2(_gnd_net_),
            .in3(N__37293),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_8_2_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_2_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIRMG61_6_LC_8_3_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIRMG61_6_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIRMG61_6_LC_8_3_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIRMG61_6_LC_8_3_0  (
            .in0(N__22438),
            .in1(N__31679),
            .in2(N__29102),
            .in3(N__30981),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNICIK32_6_LC_8_3_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNICIK32_6_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNICIK32_6_LC_8_3_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNICIK32_6_LC_8_3_1  (
            .in0(N__31681),
            .in1(N__24572),
            .in2(N__22424),
            .in3(N__24548),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNICIK32_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA8UM4_6_LC_8_3_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA8UM4_6_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA8UM4_6_LC_8_3_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA8UM4_6_LC_8_3_2  (
            .in0(N__22625),
            .in1(N__27384),
            .in2(N__22421),
            .in3(N__27628),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFJCI8_6_LC_8_3_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFJCI8_6_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFJCI8_6_LC_8_3_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFJCI8_6_LC_8_3_3  (
            .in0(N__27385),
            .in1(N__24362),
            .in2(N__22418),
            .in3(N__22598),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFJCI8_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI5T541_6_LC_8_3_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI5T541_6_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI5T541_6_LC_8_3_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI5T541_6_LC_8_3_4  (
            .in0(N__24866),
            .in1(N__31677),
            .in2(N__24890),
            .in3(N__30980),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI0VUU1_6_LC_8_3_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI0VUU1_6_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI0VUU1_6_LC_8_3_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI0VUU1_6_LC_8_3_5  (
            .in0(N__31678),
            .in1(N__22913),
            .in2(N__22628),
            .in3(N__22897),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI0VUU1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIQCIQ1_6_LC_8_3_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIQCIQ1_6_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIQCIQ1_6_LC_8_3_6 .LUT_INIT=16'b1101010110010001;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIQCIQ1_6_LC_8_3_6  (
            .in0(N__23846),
            .in1(N__31680),
            .in2(N__22619),
            .in3(N__22591),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIQCIQ1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__0_LC_8_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__0_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__0_LC_8_4_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__0_LC_8_4_0  (
            .in0(N__34799),
            .in1(N__36666),
            .in2(N__32350),
            .in3(N__32092),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33671),
            .ce(N__27774),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__1_LC_8_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__1_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__1_LC_8_4_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__1_LC_8_4_1  (
            .in0(N__36662),
            .in1(N__39596),
            .in2(N__39282),
            .in3(N__34803),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33671),
            .ce(N__27774),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__3_LC_8_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__3_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__3_LC_8_4_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__3_LC_8_4_3  (
            .in0(N__36663),
            .in1(N__34801),
            .in2(N__38188),
            .in3(N__37793),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33671),
            .ce(N__27774),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__4_LC_8_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__4_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__4_LC_8_4_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__4_LC_8_4_4  (
            .in0(N__34800),
            .in1(N__36667),
            .in2(N__35229),
            .in3(N__35546),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33671),
            .ce(N__27774),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__5_LC_8_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__5_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__5_LC_8_4_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__5_LC_8_4_5  (
            .in0(N__36664),
            .in1(N__34802),
            .in2(N__30471),
            .in3(N__30145),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33671),
            .ce(N__27774),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_5_LC_8_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_5_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_5_LC_8_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_5_LC_8_4_6  (
            .in0(N__22663),
            .in1(N__24424),
            .in2(_gnd_net_),
            .in3(N__37254),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__6_LC_8_4_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__6_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__6_LC_8_4_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__6_LC_8_4_7  (
            .in0(N__36665),
            .in1(N__29743),
            .in2(N__29370),
            .in3(N__34804),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33671),
            .ce(N__27774),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI1L181_5_LC_8_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI1L181_5_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI1L181_5_LC_8_5_0 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI1L181_5_LC_8_5_0  (
            .in0(N__28037),
            .in1(N__30837),
            .in2(N__31733),
            .in3(N__28216),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_5_LC_8_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_5_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_5_LC_8_5_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_5_LC_8_5_1  (
            .in0(N__37213),
            .in1(_gnd_net_),
            .in2(N__28217),
            .in3(N__28036),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_5_LC_8_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_5_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_5_LC_8_5_2 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_5_LC_8_5_2  (
            .in0(N__22682),
            .in1(N__28575),
            .in2(N__22709),
            .in3(N__28925),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_5_LC_8_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_5_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_5_LC_8_5_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_5_LC_8_5_3  (
            .in0(N__28576),
            .in1(N__22706),
            .in2(N__22700),
            .in3(N__22676),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_5_LC_8_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_5_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_5_LC_8_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_5_LC_8_5_4  (
            .in0(N__26443),
            .in1(N__29071),
            .in2(_gnd_net_),
            .in3(N__37211),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_5_LC_8_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_5_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_5_LC_8_5_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_5_LC_8_5_5  (
            .in0(N__37212),
            .in1(_gnd_net_),
            .in2(N__24353),
            .in3(N__26050),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI9LI91_5_LC_8_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI9LI91_5_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI9LI91_5_LC_8_5_6 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI9LI91_5_LC_8_5_6  (
            .in0(N__26051),
            .in1(N__24352),
            .in2(N__31732),
            .in3(N__30836),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIM8IQ1_5_LC_8_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIM8IQ1_5_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIM8IQ1_5_LC_8_5_7 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIM8IQ1_5_LC_8_5_7  (
            .in0(N__24425),
            .in1(N__31663),
            .in2(N__22670),
            .in3(N__22667),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIPKG61_5_LC_8_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIPKG61_5_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIPKG61_5_LC_8_6_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIPKG61_5_LC_8_6_0  (
            .in0(N__22652),
            .in1(N__31539),
            .in2(N__29816),
            .in3(N__30910),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI8EK32_5_LC_8_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI8EK32_5_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI8EK32_5_LC_8_6_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI8EK32_5_LC_8_6_1  (
            .in0(N__31541),
            .in1(N__23339),
            .in2(N__22631),
            .in3(N__23894),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_243_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI20UM4_5_LC_8_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI20UM4_5_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI20UM4_5_LC_8_6_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI20UM4_5_LC_8_6_2  (
            .in0(N__22730),
            .in1(N__27320),
            .in2(N__22808),
            .in3(N__27632),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV2CI8_5_LC_8_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV2CI8_5_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV2CI8_5_LC_8_6_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV2CI8_5_LC_8_6_3  (
            .in0(N__27321),
            .in1(N__22805),
            .in2(N__22793),
            .in3(N__22715),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI3R541_5_LC_8_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI3R541_5_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI3R541_5_LC_8_6_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNI3R541_5_LC_8_6_4  (
            .in0(N__22772),
            .in1(N__31537),
            .in2(N__24941),
            .in3(N__30909),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNISQUU1_5_LC_8_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNISQUU1_5_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNISQUU1_5_LC_8_6_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNISQUU1_5_LC_8_6_5  (
            .in0(N__31538),
            .in1(N__22949),
            .in2(N__22751),
            .in3(N__22748),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIOEMM1_5_LC_8_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIOEMM1_5_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIOEMM1_5_LC_8_6_6 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIOEMM1_5_LC_8_6_6  (
            .in0(N__26444),
            .in1(N__29075),
            .in2(N__22724),
            .in3(N__31540),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__0_LC_8_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__0_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__0_LC_8_7_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__0_LC_8_7_0  (
            .in0(N__34633),
            .in1(N__32398),
            .in2(N__32100),
            .in3(N__36403),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33651),
            .ce(N__22937),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__1_LC_8_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__1_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__1_LC_8_7_1 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__1_LC_8_7_1  (
            .in0(N__39595),
            .in1(N__34637),
            .in2(N__39290),
            .in3(N__36377),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33651),
            .ce(N__22937),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__2_LC_8_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__2_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__2_LC_8_7_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__2_LC_8_7_2  (
            .in0(N__34634),
            .in1(N__36404),
            .in2(N__38568),
            .in3(N__38799),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33651),
            .ce(N__22937),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__3_LC_8_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__3_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__3_LC_8_7_3 .LUT_INIT=16'b1100111000000010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__3_LC_8_7_3  (
            .in0(N__38118),
            .in1(N__34638),
            .in2(N__36605),
            .in3(N__37703),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33651),
            .ce(N__22937),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__4_LC_8_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__4_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__4_LC_8_7_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__4_LC_8_7_4  (
            .in0(N__34635),
            .in1(N__36405),
            .in2(N__35234),
            .in3(N__35472),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33651),
            .ce(N__22937),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__5_LC_8_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__5_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__5_LC_8_7_5 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__5_LC_8_7_5  (
            .in0(N__30069),
            .in1(N__34639),
            .in2(N__36606),
            .in3(N__30489),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33651),
            .ce(N__22937),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__6_LC_8_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__6_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__6_LC_8_7_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__6_LC_8_7_6  (
            .in0(N__34636),
            .in1(N__36406),
            .in2(N__29406),
            .in3(N__29722),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33651),
            .ce(N__22937),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_6_LC_8_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_6_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_6_LC_8_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_6_LC_8_7_7  (
            .in0(N__22909),
            .in1(N__22898),
            .in2(_gnd_net_),
            .in3(N__37356),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIUGIQ1_7_LC_8_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIUGIQ1_7_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIUGIQ1_7_LC_8_8_0 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIUGIQ1_7_LC_8_8_0  (
            .in0(N__22817),
            .in1(N__30566),
            .in2(N__22838),
            .in3(N__31684),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIUGIQ1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_7_LC_8_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_7_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_7_LC_8_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.alu_result_2_7_LC_8_8_1  (
            .in0(N__22868),
            .in1(N__22856),
            .in2(_gnd_net_),
            .in3(N__36143),
            .lcout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269 ),
            .ltout(\processor_zipi8.mux_outputs_from_alu_spm_input_ports_i.N_1269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__7_LC_8_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__7_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__7_LC_8_8_2 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__7_LC_8_8_2  (
            .in0(N__36144),
            .in1(N__33203),
            .in2(N__22841),
            .in3(N__34467),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33640),
            .ce(N__24409),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_7_LC_8_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_7_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_7_LC_8_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_7_LC_8_8_3  (
            .in0(N__37372),
            .in1(N__22834),
            .in2(_gnd_net_),
            .in3(N__22816),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIRRE01_4_LC_8_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIRRE01_4_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIRRE01_4_LC_8_8_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNIRRE01_4_LC_8_8_4  (
            .in0(N__25259),
            .in1(N__31682),
            .in2(N__25241),
            .in3(N__30898),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNICSGN1_4_LC_8_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNICSGN1_4_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNICSGN1_4_LC_8_8_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNICSGN1_4_LC_8_8_5  (
            .in0(N__31683),
            .in1(N__25220),
            .in2(N__23180),
            .in3(N__25196),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram6__RNICSGN1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_0_LC_8_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_0_LC_8_8_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe26_0_a2_0_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__27590),
            .in2(_gnd_net_),
            .in3(N__30899),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_0_LC_8_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_0_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_0_LC_8_8_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_awe28_0_a2_0_LC_8_8_7  (
            .in0(N__30900),
            .in1(_gnd_net_),
            .in2(N__27624),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_1211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_0_LC_8_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_0_LC_8_9_0 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_0_LC_8_9_0  (
            .in0(N__27001),
            .in1(N__23255),
            .in2(N__24815),
            .in3(N__28933),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_0_LC_8_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_0_LC_8_9_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_0_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__28556),
            .in2(N__23057),
            .in3(N__23051),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_1_0_LC_8_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_1_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_1_0_LC_8_9_2 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_1_0_LC_8_9_2  (
            .in0(N__30553),
            .in1(N__28931),
            .in2(N__32650),
            .in3(N__37441),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_0_LC_8_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_0_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_0_LC_8_9_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_ns_0_LC_8_9_3  (
            .in0(N__28932),
            .in1(N__24760),
            .in2(N__23054),
            .in3(N__31801),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_0_LC_8_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_0_LC_8_9_4 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_0_LC_8_9_4  (
            .in0(N__25635),
            .in1(N__25737),
            .in2(N__23045),
            .in3(N__23027),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_0_LC_8_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_0_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_0_LC_8_9_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_0_LC_8_9_5  (
            .in0(N__25636),
            .in1(N__24689),
            .in2(N__23021),
            .in3(N__23018),
            .lcout(\processor_zipi8.sy_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_1_0_LC_8_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_1_0_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_1_0_LC_8_9_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_ns_1_0_LC_8_9_6  (
            .in0(N__24719),
            .in1(N__28930),
            .in2(N__24832),
            .in3(N__37440),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_LC_8_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_LC_8_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_LC_8_10_0  (
            .in0(N__25061),
            .in1(N__26552),
            .in2(_gnd_net_),
            .in3(N__28558),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_1_LC_8_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_1_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_1_LC_8_10_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_1_LC_8_10_1  (
            .in0(N__23248),
            .in1(N__28999),
            .in2(N__23509),
            .in3(N__37451),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_LC_8_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_LC_8_10_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_LC_8_10_2  (
            .in0(N__29000),
            .in1(N__25882),
            .in2(N__23231),
            .in3(N__26032),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_LC_8_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_LC_8_10_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_LC_8_10_3  (
            .in0(N__28557),
            .in1(_gnd_net_),
            .in2(N__23228),
            .in3(N__25352),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_1_LC_8_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_1_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_1_LC_8_10_4 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_1_LC_8_10_4  (
            .in0(N__25638),
            .in1(N__23225),
            .in2(N__23216),
            .in3(N__25755),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_LC_8_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_LC_8_10_5 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_LC_8_10_5  (
            .in0(N__28559),
            .in1(N__32594),
            .in2(N__38909),
            .in3(N__24959),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_LC_8_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_LC_8_10_6 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_LC_8_10_6  (
            .in0(N__25639),
            .in1(N__23213),
            .in2(N__23207),
            .in3(N__23204),
            .lcout(\processor_zipi8.sy_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__0_LC_8_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__0_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__0_LC_8_11_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__0_LC_8_11_0  (
            .in0(N__34190),
            .in1(N__32362),
            .in2(N__32109),
            .in3(N__36192),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__1_LC_8_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__1_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__1_LC_8_11_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__1_LC_8_11_1  (
            .in0(N__36186),
            .in1(N__39450),
            .in2(N__39260),
            .in3(N__34196),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__2_LC_8_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__2_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__2_LC_8_11_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__2_LC_8_11_2  (
            .in0(N__34191),
            .in1(N__36190),
            .in2(N__38552),
            .in3(N__38878),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__3_LC_8_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__3_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__3_LC_8_11_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__3_LC_8_11_3  (
            .in0(N__36187),
            .in1(N__34194),
            .in2(N__38145),
            .in3(N__37661),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__4_LC_8_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__4_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__4_LC_8_11_4 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__4_LC_8_11_4  (
            .in0(N__34192),
            .in1(N__36191),
            .in2(N__35535),
            .in3(N__35123),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__5_LC_8_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__5_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__5_LC_8_11_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__5_LC_8_11_5  (
            .in0(N__36188),
            .in1(N__30439),
            .in2(N__30090),
            .in3(N__34197),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__6_LC_8_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__6_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__6_LC_8_11_6 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__6_LC_8_11_6  (
            .in0(N__34193),
            .in1(N__29393),
            .in2(N__29780),
            .in3(N__36193),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__7_LC_8_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__7_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__7_LC_8_11_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__7_LC_8_11_7  (
            .in0(N__36189),
            .in1(N__34195),
            .in2(N__33294),
            .in3(N__32792),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram23_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33664),
            .ce(N__23291),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__0_LC_8_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__0_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__0_LC_8_12_0 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__0_LC_8_12_0  (
            .in0(N__36279),
            .in1(N__34183),
            .in2(N__32437),
            .in3(N__32079),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33670),
            .ce(N__23438),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__1_LC_8_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__1_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__1_LC_8_12_1 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__1_LC_8_12_1  (
            .in0(N__39198),
            .in1(N__39535),
            .in2(N__34468),
            .in3(N__36284),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33670),
            .ce(N__23438),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__2_LC_8_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__2_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__2_LC_8_12_2 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__2_LC_8_12_2  (
            .in0(N__36280),
            .in1(N__38834),
            .in2(N__38530),
            .in3(N__34187),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33670),
            .ce(N__23438),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__3_LC_8_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__3_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__3_LC_8_12_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__3_LC_8_12_3  (
            .in0(N__34180),
            .in1(N__36282),
            .in2(N__37704),
            .in3(N__38078),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33670),
            .ce(N__23438),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__4_LC_8_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__4_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__4_LC_8_12_4 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__4_LC_8_12_4  (
            .in0(N__36281),
            .in1(N__35145),
            .in2(N__35556),
            .in3(N__34188),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33670),
            .ce(N__23438),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__5_LC_8_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__5_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__5_LC_8_12_5 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__5_LC_8_12_5  (
            .in0(N__34181),
            .in1(N__30067),
            .in2(N__36523),
            .in3(N__30440),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33670),
            .ce(N__23438),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_5_LC_8_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_5_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_5_LC_8_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_5_LC_8_12_6  (
            .in0(N__23722),
            .in1(N__23743),
            .in2(_gnd_net_),
            .in3(N__37505),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__6_LC_8_12_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__6_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__6_LC_8_12_7 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__6_LC_8_12_7  (
            .in0(N__34182),
            .in1(N__36283),
            .in2(N__29407),
            .in3(N__29764),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33670),
            .ce(N__23438),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__0_LC_8_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__0_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__0_LC_8_13_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__0_LC_8_13_0  (
            .in0(N__34818),
            .in1(N__32323),
            .in2(N__32080),
            .in3(N__36142),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33683),
            .ce(N__23570),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__1_LC_8_13_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__1_LC_8_13_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__1_LC_8_13_1  (
            .in0(N__36137),
            .in1(N__39568),
            .in2(N__39248),
            .in3(N__34823),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33683),
            .ce(N__23570),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__2_LC_8_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__2_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__2_LC_8_13_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__2_LC_8_13_2  (
            .in0(N__34819),
            .in1(N__36139),
            .in2(N__38461),
            .in3(N__38835),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33683),
            .ce(N__23570),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_2_LC_8_13_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_2_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_2_LC_8_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_2_LC_8_13_3  (
            .in0(N__23386),
            .in1(N__23371),
            .in2(_gnd_net_),
            .in3(N__37488),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__3_LC_8_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__3_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__3_LC_8_13_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__3_LC_8_13_4  (
            .in0(N__34820),
            .in1(N__36140),
            .in2(N__37668),
            .in3(N__38079),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33683),
            .ce(N__23570),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_3_LC_8_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_3_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_3_LC_8_13_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_am_3_LC_8_13_5  (
            .in0(N__23611),
            .in1(_gnd_net_),
            .in2(N__23596),
            .in3(N__37489),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_am_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__4_LC_8_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__4_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__4_LC_8_13_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__4_LC_8_13_6  (
            .in0(N__34821),
            .in1(N__36141),
            .in2(N__35204),
            .in3(N__35521),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33683),
            .ce(N__23570),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__5_LC_8_13_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__5_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__5_LC_8_13_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram4__5_LC_8_13_7  (
            .in0(N__36138),
            .in1(N__34822),
            .in2(N__30491),
            .in3(N__30115),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33683),
            .ce(N__23570),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__0_LC_8_14_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__0_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__0_LC_8_14_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__0_LC_8_14_0  (
            .in0(N__34810),
            .in1(N__35880),
            .in2(N__32316),
            .in3(N__31958),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__1_LC_8_14_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__1_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__1_LC_8_14_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__1_LC_8_14_1  (
            .in0(N__35876),
            .in1(N__34814),
            .in2(N__39643),
            .in3(N__39240),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__2_LC_8_14_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__2_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__2_LC_8_14_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__2_LC_8_14_2  (
            .in0(N__34811),
            .in1(N__35881),
            .in2(N__38517),
            .in3(N__38836),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__3_LC_8_14_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__3_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__3_LC_8_14_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__3_LC_8_14_3  (
            .in0(N__35877),
            .in1(N__34815),
            .in2(N__38146),
            .in3(N__37654),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__4_LC_8_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__4_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__4_LC_8_14_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__4_LC_8_14_4  (
            .in0(N__34812),
            .in1(N__35882),
            .in2(N__35231),
            .in3(N__35523),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__5_LC_8_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__5_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__5_LC_8_14_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__5_LC_8_14_5  (
            .in0(N__35878),
            .in1(N__34816),
            .in2(N__30509),
            .in3(N__30116),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__6_LC_8_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__6_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__6_LC_8_14_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__6_LC_8_14_6  (
            .in0(N__34813),
            .in1(N__35883),
            .in2(N__29408),
            .in3(N__29781),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__7_LC_8_14_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__7_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__7_LC_8_14_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram1__7_LC_8_14_7  (
            .in0(N__35879),
            .in1(N__34817),
            .in2(N__33335),
            .in3(N__32793),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33691),
            .ce(N__23762),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNITTE01_5_LC_8_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNITTE01_5_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNITTE01_5_LC_8_15_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram5__RNITTE01_5_LC_8_15_0  (
            .in0(N__23747),
            .in1(N__31612),
            .in2(N__23732),
            .in3(N__30982),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_6_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIG0HN1_5_LC_8_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIG0HN1_5_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIG0HN1_5_LC_8_15_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram6__RNIG0HN1_5_LC_8_15_1  (
            .in0(N__31613),
            .in1(N__23711),
            .in2(N__23693),
            .in3(N__23690),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNILTTE1_5_LC_8_15_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNILTTE1_5_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNILTTE1_5_LC_8_15_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNILTTE1_5_LC_8_15_2  (
            .in0(N__25048),
            .in1(N__31614),
            .in2(N__25033),
            .in3(N__30983),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI00F42_5_LC_8_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI00F42_5_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI00F42_5_LC_8_15_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNI00F42_5_LC_8_15_3  (
            .in0(N__31615),
            .in1(N__26126),
            .in2(N__23675),
            .in3(N__26114),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIENAG4_5_LC_8_15_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIENAG4_5_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIENAG4_5_LC_8_15_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__RNIENAG4_5_LC_8_15_4  (
            .in0(N__23672),
            .in1(N__27285),
            .in2(N__23666),
            .in3(N__27630),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_15_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_3_LC_8_15_5 .C_ON=1'b0;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_3_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.x12_bit_program_address_generator_i.return_vector_3_LC_8_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \processor_zipi8.x12_bit_program_address_generator_i.return_vector_3_LC_8_15_5  (
            .in0(N__23648),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\processor_zipi8.x12_bit_program_address_generator_i.return_vectorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33700),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.decode4_strobes_enables_i.un29_flag_enable_type_0_LC_8_15_6 .C_ON=1'b0;
    defparam \processor_zipi8.decode4_strobes_enables_i.un29_flag_enable_type_0_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.decode4_strobes_enables_i.un29_flag_enable_type_0_LC_8_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \processor_zipi8.decode4_strobes_enables_i.un29_flag_enable_type_0_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__24337),
            .in2(_gnd_net_),
            .in3(N__24111),
            .lcout(\processor_zipi8.un28_carry_flag_value_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__4_LC_8_16_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__4_LC_8_16_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__4_LC_8_16_4 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__4_LC_8_16_4  (
            .in0(N__36315),
            .in1(N__34189),
            .in2(N__35567),
            .in3(N__35203),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33704),
            .ce(N__25958),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__5_LC_9_2_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__5_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__5_LC_9_2_0 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__5_LC_9_2_0  (
            .in0(N__34881),
            .in1(N__36659),
            .in2(N__30155),
            .in3(N__30493),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33703),
            .ce(N__33385),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__6_LC_9_2_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__6_LC_9_2_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__6_LC_9_2_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__6_LC_9_2_1  (
            .in0(N__36658),
            .in1(N__29771),
            .in2(N__29446),
            .in3(N__34883),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33703),
            .ce(N__33385),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__7_LC_9_2_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__7_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__7_LC_9_2_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__7_LC_9_2_2  (
            .in0(N__34882),
            .in1(N__36660),
            .in2(N__33011),
            .in3(N__33339),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33703),
            .ce(N__33385),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIBNI91_6_LC_9_3_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIBNI91_6_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIBNI91_6_LC_9_3_0 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIBNI91_6_LC_9_3_0  (
            .in0(N__31674),
            .in1(N__26315),
            .in2(N__24449),
            .in3(N__30845),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_6_LC_9_3_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_6_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_6_LC_9_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_6_LC_9_3_1  (
            .in0(N__37136),
            .in1(N__28198),
            .in2(_gnd_net_),
            .in3(N__28018),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_6_LC_9_3_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_6_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_6_LC_9_3_2 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_6_LC_9_3_2  (
            .in0(N__24377),
            .in1(N__28640),
            .in2(N__23840),
            .in3(N__28973),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_6_LC_9_3_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_6_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_6_LC_9_3_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_6_LC_9_3_3  (
            .in0(N__28641),
            .in1(N__23837),
            .in2(N__23831),
            .in3(N__24371),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_6_LC_9_3_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_6_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_6_LC_9_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_6_LC_9_3_4  (
            .in0(N__26419),
            .in1(N__29053),
            .in2(_gnd_net_),
            .in3(N__37134),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_6_LC_9_3_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_6_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_6_LC_9_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_6_LC_9_3_5  (
            .in0(N__37135),
            .in1(N__26314),
            .in2(_gnd_net_),
            .in3(N__24445),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI3N181_6_LC_9_3_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI3N181_6_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI3N181_6_LC_9_3_6 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI3N181_6_LC_9_3_6  (
            .in0(N__31675),
            .in1(N__28199),
            .in2(N__28022),
            .in3(N__30846),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNISIMM1_6_LC_9_3_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNISIMM1_6_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNISIMM1_6_LC_9_3_7 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNISIMM1_6_LC_9_3_7  (
            .in0(N__29054),
            .in1(N__26420),
            .in2(N__24365),
            .in3(N__31676),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNISIMM1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__0_LC_9_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__0_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__0_LC_9_4_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__0_LC_9_4_0  (
            .in0(N__34842),
            .in1(N__36612),
            .in2(N__32351),
            .in3(N__32093),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__1_LC_9_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__1_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__1_LC_9_4_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__1_LC_9_4_1  (
            .in0(N__36608),
            .in1(N__39630),
            .in2(N__39283),
            .in3(N__34851),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__2_LC_9_4_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__2_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__2_LC_9_4_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__2_LC_9_4_2  (
            .in0(N__34843),
            .in1(N__36613),
            .in2(N__38567),
            .in3(N__38820),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__3_LC_9_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__3_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__3_LC_9_4_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__3_LC_9_4_3  (
            .in0(N__36609),
            .in1(N__34845),
            .in2(N__38189),
            .in3(N__37754),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__4_LC_9_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__4_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__4_LC_9_4_4 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__4_LC_9_4_4  (
            .in0(N__35228),
            .in1(N__35494),
            .in2(N__34880),
            .in3(N__36849),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__5_LC_9_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__5_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__5_LC_9_4_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__5_LC_9_4_5  (
            .in0(N__36610),
            .in1(N__34846),
            .in2(N__30472),
            .in3(N__30144),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__6_LC_9_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__6_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__6_LC_9_4_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__6_LC_9_4_6  (
            .in0(N__34844),
            .in1(N__36614),
            .in2(N__29369),
            .in3(N__29744),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__7_LC_9_4_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__7_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__7_LC_9_4_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__7_LC_9_4_7  (
            .in0(N__36611),
            .in1(N__33338),
            .in2(N__33028),
            .in3(N__34850),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33685),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__0_LC_9_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__0_LC_9_5_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__0_LC_9_5_0  (
            .in0(N__34618),
            .in1(N__36796),
            .in2(N__32439),
            .in3(N__32121),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33672),
            .ce(N__24408),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_0_LC_9_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_0_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_0_LC_9_5_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_0_LC_9_5_1  (
            .in0(N__24631),
            .in1(N__24652),
            .in2(_gnd_net_),
            .in3(N__37216),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__1_LC_9_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__1_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__1_LC_9_5_2 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__1_LC_9_5_2  (
            .in0(N__34619),
            .in1(N__39631),
            .in2(N__39229),
            .in3(N__36799),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33672),
            .ce(N__24408),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__2_LC_9_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__2_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__2_LC_9_5_3 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__2_LC_9_5_3  (
            .in0(N__36794),
            .in1(N__38533),
            .in2(N__38891),
            .in3(N__34624),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33672),
            .ce(N__24408),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__3_LC_9_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__3_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__3_LC_9_5_4 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__3_LC_9_5_4  (
            .in0(N__34620),
            .in1(N__36797),
            .in2(N__38187),
            .in3(N__37753),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33672),
            .ce(N__24408),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_3_LC_9_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_3_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_3_LC_9_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_3_LC_9_5_5  (
            .in0(N__26383),
            .in1(N__26365),
            .in2(_gnd_net_),
            .in3(N__37217),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__4_LC_9_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__4_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__4_LC_9_5_6 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__4_LC_9_5_6  (
            .in0(N__35093),
            .in1(N__36798),
            .in2(N__34795),
            .in3(N__35547),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33672),
            .ce(N__24408),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__5_LC_9_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__5_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__5_LC_9_5_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__5_LC_9_5_7  (
            .in0(N__36795),
            .in1(N__30448),
            .in2(N__30121),
            .in3(N__34625),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram30_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33672),
            .ce(N__24408),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_6_LC_9_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_6_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_6_LC_9_6_0 .LUT_INIT=16'b1101100001010101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_6_LC_9_6_0  (
            .in0(N__24455),
            .in1(N__24620),
            .in2(N__24530),
            .in3(N__28442),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_4_LC_9_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_4_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_4_LC_9_6_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_4_LC_9_6_1  (
            .in0(N__28060),
            .in1(N__28780),
            .in2(N__28240),
            .in3(N__37076),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_4_LC_9_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_4_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_4_LC_9_6_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_4_LC_9_6_2  (
            .in0(N__28781),
            .in1(N__26690),
            .in2(N__24596),
            .in3(N__28091),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_4_LC_9_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_4_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_4_LC_9_6_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_4_LC_9_6_3  (
            .in0(N__28440),
            .in1(_gnd_net_),
            .in2(N__24593),
            .in3(N__24467),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_6_LC_9_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_6_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_6_LC_9_6_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_6_LC_9_6_4  (
            .in0(N__37077),
            .in1(_gnd_net_),
            .in2(N__24571),
            .in3(N__24547),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_4_LC_9_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_4_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_4_LC_9_6_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_4_LC_9_6_5  (
            .in0(N__24517),
            .in1(N__28778),
            .in2(N__26074),
            .in3(N__37075),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_4_LC_9_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_4_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_4_LC_9_6_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_4_LC_9_6_6  (
            .in0(N__28779),
            .in1(N__24500),
            .in2(N__24485),
            .in3(N__24478),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_6_LC_9_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_6_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_6_LC_9_6_7 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_6_LC_9_6_7  (
            .in0(N__28441),
            .in1(N__24845),
            .in2(N__28974),
            .in3(N__24461),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNINA181_0_LC_9_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNINA181_0_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNINA181_0_LC_9_7_0 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNINA181_0_LC_9_7_0  (
            .in0(N__27749),
            .in1(N__31384),
            .in2(N__30843),
            .in3(N__27988),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_0_LC_9_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_0_LC_9_7_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_0_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__27748),
            .in2(N__27989),
            .in3(N__37089),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_0_LC_9_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_0_LC_9_7_2 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_0_LC_9_7_2  (
            .in0(N__28425),
            .in1(N__24680),
            .in2(N__24704),
            .in3(N__28774),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_0_LC_9_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_0_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_0_LC_9_7_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_0_LC_9_7_3  (
            .in0(N__24701),
            .in1(N__24674),
            .in2(N__24692),
            .in3(N__28426),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_0_LC_9_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_0_LC_9_7_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_0_LC_9_7_4  (
            .in0(N__28159),
            .in1(_gnd_net_),
            .in2(N__37245),
            .in3(N__26458),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_0_LC_9_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_0_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_0_LC_9_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_0_LC_9_7_5  (
            .in0(N__24667),
            .in1(N__26089),
            .in2(_gnd_net_),
            .in3(N__37088),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIVAI91_0_LC_9_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIVAI91_0_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIVAI91_0_LC_9_7_6 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIVAI91_0_LC_9_7_6  (
            .in0(N__26090),
            .in1(N__31385),
            .in2(N__30844),
            .in3(N__24668),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI2KHQ1_0_LC_9_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI2KHQ1_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI2KHQ1_0_LC_9_7_7 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI2KHQ1_0_LC_9_7_7  (
            .in0(N__31386),
            .in1(N__24656),
            .in2(N__24641),
            .in3(N__24638),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNI2KHQ1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIPG541_0_LC_9_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIPG541_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIPG541_0_LC_9_8_0 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIPG541_0_LC_9_8_0  (
            .in0(N__24718),
            .in1(N__31279),
            .in2(N__24836),
            .in3(N__30693),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI86UU1_0_LC_9_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI86UU1_0_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI86UU1_0_LC_9_8_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI86UU1_0_LC_9_8_1  (
            .in0(N__31280),
            .in1(N__24808),
            .in2(N__24794),
            .in3(N__27002),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNI86UU1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQMSM4_0_LC_9_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQMSM4_0_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQMSM4_0_LC_9_8_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIQMSM4_0_LC_9_8_2  (
            .in0(N__27550),
            .in1(N__27251),
            .in2(N__24791),
            .in3(N__24740),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFG9I8_0_LC_9_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFG9I8_0_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFG9I8_0_LC_9_8_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFG9I8_0_LC_9_8_3  (
            .in0(N__27252),
            .in1(N__24788),
            .in2(N__24782),
            .in3(N__24725),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFG9I8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIFAG61_0_LC_9_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIFAG61_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIFAG61_0_LC_9_8_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIFAG61_0_LC_9_8_4  (
            .in0(N__30557),
            .in1(N__31277),
            .in2(N__32651),
            .in3(N__30692),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIKPJ32_0_LC_9_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIKPJ32_0_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIKPJ32_0_LC_9_8_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIKPJ32_0_LC_9_8_5  (
            .in0(N__31278),
            .in1(N__24764),
            .in2(N__24743),
            .in3(N__31805),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIKPJ32_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI4QLM1_0_LC_9_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI4QLM1_0_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI4QLM1_0_LC_9_8_6 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI4QLM1_0_LC_9_8_6  (
            .in0(N__26462),
            .in1(N__28163),
            .in2(N__31536),
            .in3(N__24734),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI4QLM1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__0_LC_9_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__0_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__0_LC_9_9_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__0_LC_9_9_0  (
            .in0(N__34907),
            .in1(N__32349),
            .in2(N__32119),
            .in3(N__35988),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33656),
            .ce(N__24916),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__1_LC_9_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__1_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__1_LC_9_9_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__1_LC_9_9_1  (
            .in0(N__35985),
            .in1(N__34911),
            .in2(N__39619),
            .in3(N__39258),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33656),
            .ce(N__24916),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__2_LC_9_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__2_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__2_LC_9_9_2 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__2_LC_9_9_2  (
            .in0(N__34908),
            .in1(N__38550),
            .in2(N__36194),
            .in3(N__38867),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33656),
            .ce(N__24916),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__3_LC_9_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__3_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__3_LC_9_9_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__3_LC_9_9_3  (
            .in0(N__35986),
            .in1(N__34912),
            .in2(N__38172),
            .in3(N__37755),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33656),
            .ce(N__24916),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__4_LC_9_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__4_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__4_LC_9_9_4 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__4_LC_9_9_4  (
            .in0(N__34909),
            .in1(N__35189),
            .in2(N__36195),
            .in3(N__35414),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33656),
            .ce(N__24916),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__5_LC_9_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__5_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__5_LC_9_9_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__5_LC_9_9_5  (
            .in0(N__35987),
            .in1(N__34913),
            .in2(N__30498),
            .in3(N__30068),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33656),
            .ce(N__24916),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__6_LC_9_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__6_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__6_LC_9_9_6 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram17__6_LC_9_9_6  (
            .in0(N__34910),
            .in1(N__29356),
            .in2(N__29643),
            .in3(N__35989),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram17_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33656),
            .ce(N__24916),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_6_LC_9_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_6_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_6_LC_9_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_6_LC_9_9_7  (
            .in0(N__37286),
            .in1(N__24877),
            .in2(_gnd_net_),
            .in3(N__24862),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__0_LC_9_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__0_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__0_LC_9_10_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__0_LC_9_10_0  (
            .in0(N__34653),
            .in1(N__32399),
            .in2(N__32111),
            .in3(N__36548),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33665),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__1_LC_9_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__1_LC_9_10_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__1_LC_9_10_1  (
            .in0(N__36544),
            .in1(N__34654),
            .in2(N__39636),
            .in3(N__39188),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33665),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_1_LC_9_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_1_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_1_LC_9_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_1_LC_9_10_2  (
            .in0(N__37411),
            .in1(N__26794),
            .in2(_gnd_net_),
            .in3(N__26812),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__2_LC_9_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__2_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__2_LC_9_10_3 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__2_LC_9_10_3  (
            .in0(N__36545),
            .in1(N__38551),
            .in2(N__38833),
            .in3(N__34657),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33665),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_2_LC_9_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_2_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_2_LC_9_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_2_LC_9_10_4  (
            .in0(N__37410),
            .in1(N__26731),
            .in2(_gnd_net_),
            .in3(N__26752),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__3_LC_9_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__3_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__3_LC_9_10_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__3_LC_9_10_5  (
            .in0(N__36546),
            .in1(N__38067),
            .in2(N__37857),
            .in3(N__34656),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33665),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__4_LC_9_10_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__4_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__4_LC_9_10_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__4_LC_9_10_7  (
            .in0(N__36547),
            .in1(N__34655),
            .in2(N__35548),
            .in3(N__35235),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram16_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33665),
            .ce(N__25087),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_LC_9_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_LC_9_11_0 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_LC_9_11_0  (
            .in0(N__26881),
            .in1(N__24971),
            .in2(N__26861),
            .in3(N__28937),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_5_LC_9_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_5_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_5_LC_9_11_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_5_LC_9_11_1  (
            .in0(N__37450),
            .in1(_gnd_net_),
            .in2(N__25055),
            .in3(N__25034),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_5_LC_9_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_5_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_5_LC_9_11_2 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_5_LC_9_11_2  (
            .in0(N__28561),
            .in1(N__26102),
            .in2(N__25013),
            .in3(N__28939),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_5_LC_9_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_5_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_5_LC_9_11_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_5_LC_9_11_3  (
            .in0(N__25010),
            .in1(N__24995),
            .in2(N__24989),
            .in3(N__28562),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_1_LC_9_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_1_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_1_LC_9_11_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_ns_1_1_LC_9_11_4  (
            .in0(N__26536),
            .in1(N__28934),
            .in2(N__26519),
            .in3(N__37448),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_1_LC_9_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_1_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_1_LC_9_11_5 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_1_LC_9_11_5  (
            .in0(N__28938),
            .in1(N__24965),
            .in2(N__26945),
            .in3(N__28560),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_1_LC_9_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_1_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_1_LC_9_11_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_1_LC_9_11_6  (
            .in0(N__25423),
            .in1(N__28935),
            .in2(N__25406),
            .in3(N__37449),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_LC_9_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_LC_9_11_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_LC_9_11_7  (
            .in0(N__28936),
            .in1(N__25390),
            .in2(N__25373),
            .in3(N__25369),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__4_LC_9_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__4_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__4_LC_9_12_1 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__4_LC_9_12_1  (
            .in0(N__34699),
            .in1(N__35190),
            .in2(N__36599),
            .in3(N__35522),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33684),
            .ce(N__25334),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_4_LC_9_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_4_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_4_LC_9_12_2 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_1_4_LC_9_12_2  (
            .in0(N__28940),
            .in1(N__25129),
            .in2(N__25148),
            .in3(N__37249),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_4_LC_9_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_4_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_4_LC_9_12_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_ns_4_LC_9_12_3  (
            .in0(N__26185),
            .in1(N__25282),
            .in2(N__25262),
            .in3(N__28941),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_ns_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_4_LC_9_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_4_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_4_LC_9_12_4 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_1_4_LC_9_12_4  (
            .in0(N__28942),
            .in1(N__25252),
            .in2(N__25237),
            .in3(N__37250),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_4_LC_9_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_4_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_4_LC_9_12_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_6_ns_4_LC_9_12_5  (
            .in0(N__25216),
            .in1(N__25195),
            .in2(N__25172),
            .in3(N__28943),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_6_ns_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_4_LC_9_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_4_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_4_LC_9_12_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_4_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__25169),
            .in2(N__25163),
            .in3(N__28639),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIJRTE1_4_LC_9_12_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIJRTE1_4_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIJRTE1_4_LC_9_12_7 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram0__RNIJRTE1_4_LC_9_12_7  (
            .in0(N__31552),
            .in1(N__25147),
            .in2(N__25133),
            .in3(N__30916),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_2_LC_9_13_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_2_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_2_LC_9_13_0 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_2_LC_9_13_0  (
            .in0(N__28637),
            .in1(N__25838),
            .in2(N__25829),
            .in3(N__25472),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_2_LC_9_13_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_2_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_2_LC_9_13_1 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_1_2_LC_9_13_1  (
            .in0(N__25658),
            .in1(N__25814),
            .in2(N__25799),
            .in3(N__25773),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_31_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_2_LC_9_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_2_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_2_LC_9_13_2 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_31_ns_2_LC_9_13_2  (
            .in0(N__26342),
            .in1(N__25454),
            .in2(N__25673),
            .in3(N__25659),
            .lcout(\processor_zipi8.sy_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_2_LC_9_13_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_2_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_2_LC_9_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_am_2_LC_9_13_4  (
            .in0(N__37409),
            .in1(N__25504),
            .in2(_gnd_net_),
            .in3(N__25493),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_am_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_2_LC_9_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_2_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_2_LC_9_13_5 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_7_ns_1_2_LC_9_13_5  (
            .in0(N__25991),
            .in1(N__28633),
            .in2(N__25475),
            .in3(N__28944),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_7_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_2_LC_9_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_2_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_2_LC_9_13_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_2_LC_9_13_6  (
            .in0(N__28945),
            .in1(N__26903),
            .in2(N__28657),
            .in3(N__25466),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_2_LC_9_13_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_2_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_2_LC_9_13_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_2_LC_9_13_7  (
            .in0(N__38204),
            .in1(N__32558),
            .in2(N__25457),
            .in3(N__28638),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__0_LC_9_14_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__0_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__0_LC_9_14_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__0_LC_9_14_0  (
            .in0(N__34805),
            .in1(N__35885),
            .in2(N__32363),
            .in3(N__31959),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33702),
            .ce(N__25957),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__1_LC_9_14_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__1_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__1_LC_9_14_1 .LUT_INIT=16'b1010101000001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__1_LC_9_14_1  (
            .in0(N__39241),
            .in1(N__39626),
            .in2(N__36098),
            .in3(N__34808),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33702),
            .ce(N__25957),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__2_LC_9_14_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__2_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__2_LC_9_14_2 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__2_LC_9_14_2  (
            .in0(N__34806),
            .in1(N__38782),
            .in2(N__36099),
            .in3(N__38425),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33702),
            .ce(N__25957),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_2_LC_9_14_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_2_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_2_LC_9_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_2_LC_9_14_3  (
            .in0(N__25849),
            .in1(N__26002),
            .in2(_gnd_net_),
            .in3(N__37478),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__3_LC_9_14_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__3_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__3_LC_9_14_4 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__3_LC_9_14_4  (
            .in0(N__34807),
            .in1(N__35886),
            .in2(N__38173),
            .in3(N__37629),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33702),
            .ce(N__25957),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_3_LC_9_14_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_3_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_3_LC_9_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_3_LC_9_14_5  (
            .in0(N__26200),
            .in1(N__25981),
            .in2(_gnd_net_),
            .in3(N__37477),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__5_LC_9_14_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__5_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__5_LC_9_14_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram2__5_LC_9_14_7  (
            .in0(N__35884),
            .in1(N__30494),
            .in2(N__30150),
            .in3(N__34809),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33702),
            .ce(N__25957),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__0_LC_9_15_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__0_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__0_LC_9_15_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__0_LC_9_15_0  (
            .in0(N__33926),
            .in1(N__36312),
            .in2(N__32364),
            .in3(N__32058),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33705),
            .ce(N__26168),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__1_LC_9_15_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__1_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__1_LC_9_15_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__1_LC_9_15_1  (
            .in0(N__36309),
            .in1(N__33929),
            .in2(N__39645),
            .in3(N__39226),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33705),
            .ce(N__26168),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__2_LC_9_15_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__2_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__2_LC_9_15_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__2_LC_9_15_2  (
            .in0(N__33927),
            .in1(N__36313),
            .in2(N__38531),
            .in3(N__38783),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33705),
            .ce(N__26168),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__3_LC_9_15_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__3_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__3_LC_9_15_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__3_LC_9_15_3  (
            .in0(N__36310),
            .in1(N__33930),
            .in2(N__38186),
            .in3(N__37705),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33705),
            .ce(N__26168),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__4_LC_9_15_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__4_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__4_LC_9_15_4 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__4_LC_9_15_4  (
            .in0(N__33928),
            .in1(N__35220),
            .in2(N__35568),
            .in3(N__36314),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33705),
            .ce(N__26168),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__5_LC_9_15_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__5_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__5_LC_9_15_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram3__5_LC_9_15_5  (
            .in0(N__36311),
            .in1(N__33931),
            .in2(N__30510),
            .in3(N__30117),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33705),
            .ce(N__26168),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_5_LC_9_15_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_5_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_5_LC_9_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_3_bm_5_LC_9_15_6  (
            .in0(N__26125),
            .in1(N__26113),
            .in2(_gnd_net_),
            .in3(N__37490),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_3_bm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__0_LC_11_4_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__0_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__0_LC_11_4_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__0_LC_11_4_0  (
            .in0(N__34610),
            .in1(N__36619),
            .in2(N__32352),
            .in3(N__32123),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__1_LC_11_4_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__1_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__1_LC_11_4_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__1_LC_11_4_1  (
            .in0(N__36615),
            .in1(N__39637),
            .in2(N__39284),
            .in3(N__34616),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__2_LC_11_4_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__2_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__2_LC_11_4_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__2_LC_11_4_2  (
            .in0(N__34611),
            .in1(N__36620),
            .in2(N__38576),
            .in3(N__38889),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__3_LC_11_4_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__3_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__3_LC_11_4_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__3_LC_11_4_3  (
            .in0(N__36616),
            .in1(N__34614),
            .in2(N__38192),
            .in3(N__37778),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__4_LC_11_4_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__4_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__4_LC_11_4_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__4_LC_11_4_4  (
            .in0(N__34612),
            .in1(N__36621),
            .in2(N__35232),
            .in3(N__35428),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__5_LC_11_4_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__5_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__5_LC_11_4_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__5_LC_11_4_5  (
            .in0(N__36617),
            .in1(N__34615),
            .in2(N__30473),
            .in3(N__30154),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__6_LC_11_4_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__6_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__6_LC_11_4_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__6_LC_11_4_6  (
            .in0(N__34613),
            .in1(N__36622),
            .in2(N__29368),
            .in3(N__29772),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__7_LC_11_4_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__7_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__7_LC_11_4_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram29__7_LC_11_4_7  (
            .in0(N__36618),
            .in1(N__33334),
            .in2(N__33001),
            .in3(N__34617),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33697),
            .ce(N__26294),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNITG181_3_LC_11_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNITG181_3_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNITG181_3_LC_11_5_0 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNITG181_3_LC_11_5_0  (
            .in0(N__28070),
            .in1(N__31515),
            .in2(N__30979),
            .in3(N__27941),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_3_LC_11_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_3_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_3_LC_11_5_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_3_LC_11_5_1  (
            .in0(N__37071),
            .in1(N__27094),
            .in2(_gnd_net_),
            .in3(N__28108),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_3_LC_11_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_3_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_3_LC_11_5_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_3_LC_11_5_2  (
            .in0(N__26246),
            .in1(N__28527),
            .in2(N__26282),
            .in3(N__28893),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_3_LC_11_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_3_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_3_LC_11_5_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_3_LC_11_5_3  (
            .in0(N__28528),
            .in1(N__26279),
            .in2(N__26270),
            .in3(N__26240),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_3_LC_11_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_3_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_3_LC_11_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_3_LC_11_5_4  (
            .in0(N__28069),
            .in1(N__27940),
            .in2(_gnd_net_),
            .in3(N__37069),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_3_LC_11_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_3_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_3_LC_11_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_3_LC_11_5_5  (
            .in0(N__37070),
            .in1(N__26215),
            .in2(_gnd_net_),
            .in3(N__26233),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI5HI91_3_LC_11_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI5HI91_3_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI5HI91_3_LC_11_5_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI5HI91_3_LC_11_5_6  (
            .in0(N__26234),
            .in1(N__31516),
            .in2(N__26219),
            .in3(N__30864),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIE0IQ1_3_LC_11_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIE0IQ1_3_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIE0IQ1_3_LC_11_5_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIE0IQ1_3_LC_11_5_7  (
            .in0(N__31517),
            .in1(N__26390),
            .in2(N__26372),
            .in3(N__26369),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIE0IQ1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_2_LC_11_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_2_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_2_LC_11_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_bm_2_LC_11_6_0  (
            .in0(N__27808),
            .in1(N__26602),
            .in2(_gnd_net_),
            .in3(N__37066),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIRE181_2_LC_11_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIRE181_2_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIRE181_2_LC_11_6_1 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIRE181_2_LC_11_6_1  (
            .in0(N__27716),
            .in1(N__31507),
            .in2(N__30943),
            .in3(N__27950),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_2_LC_11_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_2_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_2_LC_11_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_2_LC_11_6_2  (
            .in0(N__27949),
            .in1(N__27715),
            .in2(_gnd_net_),
            .in3(N__37068),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_2_LC_11_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_2_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_2_LC_11_6_3 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_2_LC_11_6_3  (
            .in0(N__28767),
            .in1(N__26327),
            .in2(N__26354),
            .in3(N__28427),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_2_LC_11_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_2_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_2_LC_11_6_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_2_LC_11_6_4  (
            .in0(N__28428),
            .in1(N__26351),
            .in2(N__26345),
            .in3(N__26321),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_2_LC_11_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_2_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_2_LC_11_6_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_2_LC_11_6_5  (
            .in0(N__37064),
            .in1(_gnd_net_),
            .in2(N__28129),
            .in3(N__26716),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_1_LC_11_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_1_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_1_LC_11_6_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_1_LC_11_6_6  (
            .in0(N__27727),
            .in1(N__28766),
            .in2(N__27967),
            .in3(N__37065),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_2_LC_11_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_2_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_2_LC_11_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_2_LC_11_6_7  (
            .in0(N__37067),
            .in1(N__26620),
            .in2(_gnd_net_),
            .in3(N__26647),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__0_LC_11_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__0_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__0_LC_11_7_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__0_LC_11_7_0  (
            .in0(N__34582),
            .in1(N__36382),
            .in2(N__32474),
            .in3(N__32088),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__1_LC_11_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__1_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__1_LC_11_7_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__1_LC_11_7_1  (
            .in0(N__36378),
            .in1(N__39608),
            .in2(N__39289),
            .in3(N__34586),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__2_LC_11_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__2_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__2_LC_11_7_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__2_LC_11_7_2  (
            .in0(N__34583),
            .in1(N__36383),
            .in2(N__38569),
            .in3(N__38800),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__3_LC_11_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__3_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__3_LC_11_7_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__3_LC_11_7_3  (
            .in0(N__36379),
            .in1(N__38136),
            .in2(N__37835),
            .in3(N__34587),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__4_LC_11_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__4_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__4_LC_11_7_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__4_LC_11_7_4  (
            .in0(N__34584),
            .in1(N__36384),
            .in2(N__35236),
            .in3(N__35498),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__5_LC_11_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__5_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__5_LC_11_7_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__5_LC_11_7_5  (
            .in0(N__36380),
            .in1(N__30477),
            .in2(N__30136),
            .in3(N__34588),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__6_LC_11_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__6_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__6_LC_11_7_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__6_LC_11_7_6  (
            .in0(N__34585),
            .in1(N__36385),
            .in2(N__29395),
            .in3(N__29708),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__7_LC_11_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__7_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__7_LC_11_7_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram27__7_LC_11_7_7  (
            .in0(N__36381),
            .in1(N__33290),
            .in2(N__32999),
            .in3(N__34589),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33666),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIVI181_4_LC_11_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIVI181_4_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIVI181_4_LC_11_8_0 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIVI181_4_LC_11_8_0  (
            .in0(N__30659),
            .in1(N__28061),
            .in2(N__28244),
            .in3(N__31341),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIKAMM1_4_LC_11_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIKAMM1_4_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIKAMM1_4_LC_11_8_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIKAMM1_4_LC_11_8_1  (
            .in0(N__31342),
            .in1(N__26689),
            .in2(N__26669),
            .in3(N__28084),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIKAMM1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIPC181_1_LC_11_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIPC181_1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIPC181_1_LC_11_8_2 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNIPC181_1_LC_11_8_2  (
            .in0(N__30656),
            .in1(N__27734),
            .in2(N__27971),
            .in3(N__31337),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI8ULM1_1_LC_11_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI8ULM1_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI8ULM1_1_LC_11_8_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI8ULM1_1_LC_11_8_3  (
            .in0(N__31338),
            .in1(N__26579),
            .in2(N__26651),
            .in3(N__28142),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI3FI91_2_LC_11_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI3FI91_2_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI3FI91_2_LC_11_8_4 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI3FI91_2_LC_11_8_4  (
            .in0(N__30658),
            .in1(N__26648),
            .in2(N__26624),
            .in3(N__31339),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIASHQ1_2_LC_11_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIASHQ1_2_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIASHQ1_2_LC_11_8_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNIASHQ1_2_LC_11_8_5  (
            .in0(N__31340),
            .in1(N__27809),
            .in2(N__26606),
            .in3(N__26603),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram30__RNIASHQ1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_LC_11_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_LC_11_8_6 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_ns_1_LC_11_8_6  (
            .in0(N__28141),
            .in1(N__26578),
            .in2(N__26564),
            .in3(N__28889),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI1DI91_1_LC_11_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI1DI91_1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI1DI91_1_LC_11_8_7 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNI1DI91_1_LC_11_8_7  (
            .in0(N__31336),
            .in1(N__26540),
            .in2(N__26515),
            .in3(N__30657),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI2VSM4_1_LC_11_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI2VSM4_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI2VSM4_1_LC_11_9_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNI2VSM4_1_LC_11_9_0  (
            .in0(N__26780),
            .in1(N__27191),
            .in2(N__26768),
            .in3(N__27540),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV0AI8_1_LC_11_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV0AI8_1_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV0AI8_1_LC_11_9_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV0AI8_1_LC_11_9_1  (
            .in0(N__27192),
            .in1(N__26489),
            .in2(N__26480),
            .in3(N__26825),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI6OHQ1_1_LC_11_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI6OHQ1_1_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI6OHQ1_1_LC_11_9_2 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram30__RNI6OHQ1_1_LC_11_9_2  (
            .in0(N__26891),
            .in1(N__26867),
            .in2(N__26860),
            .in3(N__31175),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIHCG61_1_LC_11_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIHCG61_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIHCG61_1_LC_11_9_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIHCG61_1_LC_11_9_3  (
            .in0(N__30635),
            .in1(N__32621),
            .in2(N__31305),
            .in3(N__32605),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIRI541_1_LC_11_9_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIRI541_1_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIRI541_1_LC_11_9_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIRI541_1_LC_11_9_4  (
            .in0(N__26819),
            .in1(N__31172),
            .in2(N__26801),
            .in3(N__30636),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNICAUU1_1_LC_11_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNICAUU1_1_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNICAUU1_1_LC_11_9_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNICAUU1_1_LC_11_9_5  (
            .in0(N__31173),
            .in1(N__26978),
            .in2(N__26783),
            .in3(N__26960),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIOTJ32_1_LC_11_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIOTJ32_1_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIOTJ32_1_LC_11_9_6 .LUT_INIT=16'b1101100001010101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIOTJ32_1_LC_11_9_6  (
            .in0(N__26774),
            .in1(N__38924),
            .in2(N__38948),
            .in3(N__31174),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIJEG61_2_LC_11_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIJEG61_2_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIJEG61_2_LC_11_10_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNIJEG61_2_LC_11_10_0  (
            .in0(N__32570),
            .in1(N__31217),
            .in2(N__32585),
            .in3(N__30690),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIS1K32_2_LC_11_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIS1K32_2_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIS1K32_2_LC_11_10_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNIS1K32_2_LC_11_10_1  (
            .in0(N__31219),
            .in1(N__38219),
            .in2(N__26759),
            .in3(N__38240),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNIS1K32_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNITK541_2_LC_11_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNITK541_2_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNITK541_2_LC_11_10_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNITK541_2_LC_11_10_2  (
            .in0(N__26756),
            .in1(N__31218),
            .in2(N__26741),
            .in3(N__30691),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIC2MM1_2_LC_11_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIC2MM1_2_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIC2MM1_2_LC_11_10_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIC2MM1_2_LC_11_10_3  (
            .in0(N__31221),
            .in1(N__26720),
            .in2(N__26705),
            .in3(N__28133),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIC2MM1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFHAI8_2_LC_11_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFHAI8_2_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFHAI8_2_LC_11_10_4 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIFHAI8_2_LC_11_10_4  (
            .in0(N__27059),
            .in1(N__27008),
            .in2(N__27044),
            .in3(N__27206),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIFHAI8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIGEUU1_2_LC_11_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIGEUU1_2_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIGEUU1_2_LC_11_10_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIGEUU1_2_LC_11_10_5  (
            .in0(N__31220),
            .in1(N__26933),
            .in2(N__27026),
            .in3(N__26915),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIGEUU1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA7TM4_2_LC_11_10_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA7TM4_2_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA7TM4_2_LC_11_10_6 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIA7TM4_2_LC_11_10_6  (
            .in0(N__27541),
            .in1(N__27017),
            .in2(N__27011),
            .in3(N__27205),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__0_LC_11_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__0_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__0_LC_11_11_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__0_LC_11_11_0  (
            .in0(N__34203),
            .in1(N__36185),
            .in2(N__32476),
            .in3(N__32102),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33686),
            .ce(N__27686),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__1_LC_11_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__1_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__1_LC_11_11_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__1_LC_11_11_1  (
            .in0(N__36181),
            .in1(N__34204),
            .in2(N__39542),
            .in3(N__39261),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33686),
            .ce(N__27686),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_1_LC_11_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_1_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_1_LC_11_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_1_LC_11_11_2  (
            .in0(N__26977),
            .in1(N__26956),
            .in2(_gnd_net_),
            .in3(N__37432),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__2_LC_11_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__2_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__2_LC_11_11_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__2_LC_11_11_3  (
            .in0(N__36182),
            .in1(N__38831),
            .in2(N__38570),
            .in3(N__34207),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33686),
            .ce(N__27686),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_2_LC_11_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_2_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_2_LC_11_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_2_LC_11_11_4  (
            .in0(N__26932),
            .in1(N__26914),
            .in2(_gnd_net_),
            .in3(N__37430),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__3_LC_11_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__3_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__3_LC_11_11_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__3_LC_11_11_5  (
            .in0(N__36183),
            .in1(N__34205),
            .in2(N__38182),
            .in3(N__37702),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33686),
            .ce(N__27686),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_3_LC_11_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_3_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_3_LC_11_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_bm_3_LC_11_11_6  (
            .in0(N__27928),
            .in1(N__27907),
            .in2(_gnd_net_),
            .in3(N__37431),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_bm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__4_LC_11_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__4_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__4_LC_11_11_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram18__4_LC_11_11_7  (
            .in0(N__36184),
            .in1(N__34206),
            .in2(N__35559),
            .in3(N__35170),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram18_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33686),
            .ce(N__27686),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNILGG61_3_LC_11_12_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNILGG61_3_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNILGG61_3_LC_11_12_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__RNILGG61_3_LC_11_12_0  (
            .in0(N__30798),
            .in1(N__30536),
            .in2(N__31508),
            .in3(N__32545),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_21_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI06K32_3_LC_11_12_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI06K32_3_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI06K32_3_LC_11_12_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram23__RNI06K32_3_LC_11_12_1  (
            .in0(N__37538),
            .in1(N__37517),
            .in2(N__27647),
            .in3(N__31326),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram23__RNI06K32_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIFTM4_3_LC_11_12_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIFTM4_3_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIFTM4_3_LC_11_12_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIIFTM4_3_LC_11_12_2  (
            .in0(N__27896),
            .in1(N__27186),
            .in2(N__27644),
            .in3(N__27539),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_30_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV1BI8_3_LC_11_12_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV1BI8_3_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV1BI8_3_LC_11_12_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIV1BI8_3_LC_11_12_3  (
            .in0(N__27187),
            .in1(N__27122),
            .in2(N__27113),
            .in3(N__27065),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIV1BI8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIG6MM1_3_LC_11_12_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIG6MM1_3_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIG6MM1_3_LC_11_12_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNIG6MM1_3_LC_11_12_4  (
            .in0(N__31325),
            .in1(N__27095),
            .in2(N__27077),
            .in3(N__28112),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNIG6MM1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIVM541_3_LC_11_12_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIVM541_3_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIVM541_3_LC_11_12_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram16__RNIVM541_3_LC_11_12_5  (
            .in0(N__27866),
            .in1(N__31320),
            .in2(N__27890),
            .in3(N__30797),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_18_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIKIUU1_3_LC_11_12_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIKIUU1_3_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIKIUU1_3_LC_11_12_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram19__RNIKIUU1_3_LC_11_12_6  (
            .in0(N__31321),
            .in1(N__27932),
            .in2(N__27911),
            .in3(N__27908),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram19__RNIKIUU1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_3_LC_11_13_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_3_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_3_LC_11_13_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_3_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__37438),
            .in2(N__32546),
            .in3(N__30535),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_3_LC_11_13_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_3_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_3_LC_11_13_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_18_am_3_LC_11_13_5  (
            .in0(N__27886),
            .in1(N__37439),
            .in2(_gnd_net_),
            .in3(N__27865),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_18_am_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_3_LC_11_13_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_3_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_3_LC_11_13_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_1_3_LC_11_13_6  (
            .in0(N__27842),
            .in1(N__28613),
            .in2(N__27833),
            .in3(N__28969),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_3_LC_11_13_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_3_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_3_LC_11_13_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_22_ns_3_LC_11_13_7  (
            .in0(N__28614),
            .in1(N__36866),
            .in2(N__27830),
            .in3(N__27827),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_22_ns_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__2_LC_11_14_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__2_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__2_LC_11_14_6 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram31__2_LC_11_14_6  (
            .in0(N__34726),
            .in1(N__38505),
            .in2(N__36100),
            .in3(N__38832),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram31_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33710),
            .ce(N__27788),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__0_LC_12_5_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__0_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__0_LC_12_5_0 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__0_LC_12_5_0  (
            .in0(N__32120),
            .in1(N__32438),
            .in2(N__34794),
            .in3(N__36847),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__1_LC_12_5_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__1_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__1_LC_12_5_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__1_LC_12_5_1  (
            .in0(N__36840),
            .in1(N__34600),
            .in2(N__39646),
            .in3(N__39263),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__2_LC_12_5_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__2_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__2_LC_12_5_2 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__2_LC_12_5_2  (
            .in0(N__38882),
            .in1(N__36844),
            .in2(N__34793),
            .in3(N__38574),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__3_LC_12_5_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__3_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__3_LC_12_5_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__3_LC_12_5_3  (
            .in0(N__36841),
            .in1(N__34601),
            .in2(N__38191),
            .in3(N__37810),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__4_LC_12_5_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__4_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__4_LC_12_5_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__4_LC_12_5_4  (
            .in0(N__34598),
            .in1(N__36845),
            .in2(N__35169),
            .in3(N__35545),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__5_LC_12_5_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__5_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__5_LC_12_5_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__5_LC_12_5_5  (
            .in0(N__36842),
            .in1(N__34602),
            .in2(N__30514),
            .in3(N__30147),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__6_LC_12_5_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__6_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__6_LC_12_5_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__6_LC_12_5_6  (
            .in0(N__34599),
            .in1(N__36846),
            .in2(N__29437),
            .in3(N__29751),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__7_LC_12_5_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__7_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__7_LC_12_5_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__7_LC_12_5_7  (
            .in0(N__36843),
            .in1(N__33333),
            .in2(N__32960),
            .in3(N__34609),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram24_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33699),
            .ce(N__28004),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__0_LC_12_6_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__0_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__0_LC_12_6_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__0_LC_12_6_0  (
            .in0(N__34590),
            .in1(N__36740),
            .in2(N__32475),
            .in3(N__32122),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__1_LC_12_6_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__1_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__1_LC_12_6_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__1_LC_12_6_1  (
            .in0(N__36736),
            .in1(N__34594),
            .in2(N__39638),
            .in3(N__39243),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__2_LC_12_6_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__2_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__2_LC_12_6_2 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__2_LC_12_6_2  (
            .in0(N__34591),
            .in1(N__36741),
            .in2(N__38888),
            .in3(N__38575),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__3_LC_12_6_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__3_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__3_LC_12_6_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__3_LC_12_6_3  (
            .in0(N__36737),
            .in1(N__34595),
            .in2(N__38190),
            .in3(N__37756),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__4_LC_12_6_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__4_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__4_LC_12_6_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__4_LC_12_6_4  (
            .in0(N__34592),
            .in1(N__36742),
            .in2(N__35233),
            .in3(N__35485),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__5_LC_12_6_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__5_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__5_LC_12_6_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__5_LC_12_6_5  (
            .in0(N__36738),
            .in1(N__34596),
            .in2(N__30518),
            .in3(N__30148),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__6_LC_12_6_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__6_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__6_LC_12_6_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__6_LC_12_6_6  (
            .in0(N__34593),
            .in1(N__36743),
            .in2(N__29394),
            .in3(N__29710),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__7_LC_12_6_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__7_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__7_LC_12_6_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram25__7_LC_12_6_7  (
            .in0(N__36739),
            .in1(N__34597),
            .in2(N__33336),
            .in3(N__32944),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram25_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33688),
            .ce(N__28181),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__0_LC_12_7_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__0_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__0_LC_12_7_0 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__0_LC_12_7_0  (
            .in0(N__34884),
            .in1(N__32461),
            .in2(N__36851),
            .in3(N__32087),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__1_LC_12_7_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__1_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__1_LC_12_7_1 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__1_LC_12_7_1  (
            .in0(N__34885),
            .in1(N__39609),
            .in2(N__39285),
            .in3(N__36830),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__2_LC_12_7_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__2_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__2_LC_12_7_2 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__2_LC_12_7_2  (
            .in0(N__38541),
            .in1(N__34890),
            .in2(N__36852),
            .in3(N__38801),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__3_LC_12_7_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__3_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__3_LC_12_7_3 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__3_LC_12_7_3  (
            .in0(N__34886),
            .in1(N__36819),
            .in2(N__38181),
            .in3(N__37823),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__4_LC_12_7_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__4_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__4_LC_12_7_4 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__4_LC_12_7_4  (
            .in0(N__36818),
            .in1(N__35221),
            .in2(N__35558),
            .in3(N__34891),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__5_LC_12_7_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__5_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__5_LC_12_7_5 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__5_LC_12_7_5  (
            .in0(N__34887),
            .in1(N__30481),
            .in2(N__30135),
            .in3(N__36829),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__6_LC_12_7_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__6_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__6_LC_12_7_6 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__6_LC_12_7_6  (
            .in0(N__29398),
            .in1(N__34889),
            .in2(N__36853),
            .in3(N__29709),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__7_LC_12_7_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__7_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__7_LC_12_7_7 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__7_LC_12_7_7  (
            .in0(N__34888),
            .in1(N__32872),
            .in2(N__33317),
            .in3(N__36831),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram26_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33677),
            .ce(N__29036),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_7_LC_12_8_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_7_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_7_LC_12_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_28_am_7_LC_12_8_0  (
            .in0(N__31039),
            .in1(N__31060),
            .in2(_gnd_net_),
            .in3(N__37252),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_28_am_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_7_LC_12_8_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_7_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_7_LC_12_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_am_7_LC_12_8_1  (
            .in0(N__37253),
            .in1(N__28291),
            .in2(_gnd_net_),
            .in3(N__28273),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_am_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_7_LC_12_8_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_7_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_7_LC_12_8_2 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_1_7_LC_12_8_2  (
            .in0(N__31757),
            .in1(N__28615),
            .in2(N__29018),
            .in3(N__29003),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_7_LC_12_8_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_7_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_7_LC_12_8_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_29_ns_7_LC_12_8_3  (
            .in0(N__28616),
            .in1(N__28331),
            .in2(N__28319),
            .in3(N__28316),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_29_ns_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI5P181_7_LC_12_8_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI5P181_7_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI5P181_7_LC_12_8_4 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram24__RNI5P181_7_LC_12_8_4  (
            .in0(N__30860),
            .in1(N__28292),
            .in2(N__28277),
            .in3(N__31691),
            .lcout(),
            .ltout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_25_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI0NMM1_7_LC_12_8_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI0NMM1_7_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI0NMM1_7_LC_12_8_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram26__RNI0NMM1_7_LC_12_8_5  (
            .in0(N__31692),
            .in1(N__31768),
            .in2(N__28262),
            .in3(N__31778),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_ram26__RNI0NMM1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_7_LC_12_8_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_7_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_7_LC_12_8_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_25_bm_7_LC_12_8_6  (
            .in0(N__31777),
            .in1(_gnd_net_),
            .in2(N__31769),
            .in3(N__37251),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_25_bm_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIDPI91_7_LC_12_8_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIDPI91_7_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIDPI91_7_LC_12_8_7 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram28__RNIDPI91_7_LC_12_8_7  (
            .in0(N__31690),
            .in1(N__31061),
            .in2(N__31043),
            .in3(N__30859),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ramout_28_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__0_LC_12_9_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__0_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__0_LC_12_9_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__0_LC_12_9_0  (
            .in0(N__34832),
            .in1(N__35994),
            .in2(N__32458),
            .in3(N__32110),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33678),
            .ce(N__32684),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__1_LC_12_9_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__1_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__1_LC_12_9_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__1_LC_12_9_1  (
            .in0(N__35990),
            .in1(N__34835),
            .in2(N__39642),
            .in3(N__39177),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33678),
            .ce(N__32684),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__2_LC_12_9_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__2_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__2_LC_12_9_2 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__2_LC_12_9_2  (
            .in0(N__34833),
            .in1(N__38887),
            .in2(N__36854),
            .in3(N__38565),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33678),
            .ce(N__32684),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__3_LC_12_9_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__3_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__3_LC_12_9_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__3_LC_12_9_3  (
            .in0(N__35991),
            .in1(N__38137),
            .in2(N__37840),
            .in3(N__34838),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33678),
            .ce(N__32684),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__5_LC_12_9_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__5_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__5_LC_12_9_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__5_LC_12_9_5  (
            .in0(N__35992),
            .in1(N__34836),
            .in2(N__30507),
            .in3(N__30149),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33678),
            .ce(N__32684),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__6_LC_12_9_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__6_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__6_LC_12_9_6 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__6_LC_12_9_6  (
            .in0(N__34834),
            .in1(N__35995),
            .in2(N__29768),
            .in3(N__29438),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33678),
            .ce(N__32684),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__7_LC_12_9_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__7_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__7_LC_12_9_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram21__7_LC_12_9_7  (
            .in0(N__35993),
            .in1(N__34837),
            .in2(N__33337),
            .in3(N__33000),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram21_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33678),
            .ce(N__32684),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__0_LC_12_10_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__0_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__0_LC_12_10_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__0_LC_12_10_0  (
            .in0(N__34701),
            .in1(N__36836),
            .in2(N__32459),
            .in3(N__32115),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33687),
            .ce(N__32507),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__1_LC_12_10_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__1_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__1_LC_12_10_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__1_LC_12_10_1  (
            .in0(N__36832),
            .in1(N__34702),
            .in2(N__39647),
            .in3(N__39242),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33687),
            .ce(N__32507),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_1_LC_12_10_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_1_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_1_LC_12_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_1_LC_12_10_2  (
            .in0(N__32620),
            .in1(N__32606),
            .in2(_gnd_net_),
            .in3(N__37397),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__2_LC_12_10_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__2_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__2_LC_12_10_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__2_LC_12_10_3  (
            .in0(N__36833),
            .in1(N__34703),
            .in2(N__38843),
            .in3(N__38566),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33687),
            .ce(N__32507),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_2_LC_12_10_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_2_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_2_LC_12_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_am_2_LC_12_10_4  (
            .in0(N__32581),
            .in1(N__32569),
            .in2(_gnd_net_),
            .in3(N__37396),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_am_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__3_LC_12_10_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__3_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__3_LC_12_10_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__3_LC_12_10_5  (
            .in0(N__36834),
            .in1(N__38122),
            .in2(N__37858),
            .in3(N__34831),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33687),
            .ce(N__32507),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__4_LC_12_10_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__4_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__4_LC_12_10_7 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram20__4_LC_12_10_7  (
            .in0(N__36835),
            .in1(N__34704),
            .in2(N__35557),
            .in3(N__35240),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33687),
            .ce(N__32507),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__0_LC_12_11_0 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__0_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__0_LC_12_11_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__0_LC_12_11_0  (
            .in0(N__34198),
            .in1(N__36604),
            .in2(N__32477),
            .in3(N__32101),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33698),
            .ce(N__33389),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__1_LC_12_11_1 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__1_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__1_LC_12_11_1 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__1_LC_12_11_1  (
            .in0(N__36600),
            .in1(N__34199),
            .in2(N__39543),
            .in3(N__39259),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33698),
            .ce(N__33389),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_1_LC_12_11_2 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_1_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_1_LC_12_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_1_LC_12_11_2  (
            .in0(N__38941),
            .in1(N__38920),
            .in2(_gnd_net_),
            .in3(N__37502),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__2_LC_12_11_3 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__2_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__2_LC_12_11_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__2_LC_12_11_3  (
            .in0(N__36601),
            .in1(N__34200),
            .in2(N__38890),
            .in3(N__38549),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33698),
            .ce(N__33389),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_2_LC_12_11_4 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_2_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_2_LC_12_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_2_LC_12_11_4  (
            .in0(N__38236),
            .in1(N__38215),
            .in2(_gnd_net_),
            .in3(N__37500),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__3_LC_12_11_5 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__3_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__3_LC_12_11_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__3_LC_12_11_5  (
            .in0(N__36602),
            .in1(N__34201),
            .in2(N__38183),
            .in3(N__37836),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33698),
            .ce(N__33389),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_3_LC_12_11_6 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_3_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_3_LC_12_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ram_s_rd_wr_ramout_21_bm_3_LC_12_11_6  (
            .in0(N__37534),
            .in1(N__37516),
            .in2(_gnd_net_),
            .in3(N__37501),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.sy_bank.ramout_21_bm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__4_LC_12_11_7 .C_ON=1'b0;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__4_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__4_LC_12_11_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \processor_zipi8.two_banks_of_16_gp_reg_i.sx_bank.ram_s_two_banks_of_16_gp_reg_i_sx_bank_ram_s_ram22__4_LC_12_11_7  (
            .in0(N__36603),
            .in1(N__35531),
            .in2(N__35219),
            .in3(N__34202),
            .lcout(\processor_zipi8.two_banks_of_16_gp_reg_i.ram22_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33698),
            .ce(N__33389),
            .sr(_gnd_net_));
endmodule // top
