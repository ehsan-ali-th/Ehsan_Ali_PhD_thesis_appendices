// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Jul 10 03:17:48 2019
//
// Verilog Description of module top
//

module top (CLK_3P3_MHZ, BTN1, LED1);   // src/top.vhd(34[8:11])
    input CLK_3P3_MHZ;   // src/top.vhd(36[9:20])
    input BTN1;   // src/top.vhd(37[9:13])
    output LED1;   // src/top.vhd(38[3:7])
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    wire GND_net, BTN1_c, LED1_c_0;
    wire [11:0]address;   // src/top.vhd(80[20:27])
    wire [17:0]instruction;   // src/top.vhd(81[16:27])
    
    wire bram_enable, ram_s_36_5, ram_s_36_4, ram_s_36_3, ram_s_44_1, 
        ram_s_44_0, ram_s_43_7, ram_s_43_6, ram_s_43_5, ram_s_43_4, 
        ram_s_43_3, ram_s_43_2, ram_s_43_1, ram_s_43_0;
    wire [2:1]t_state;   // src/zipi8.vhd(279[12:19])
    
    wire ram_s_32_6, internal_reset, n899, ram_s_36_6, ram_s_32_0;
    wire [11:0]register_vector;   // src/zipi8.vhd(312[12:27])
    
    wire special_bit;
    wire [7:0]sx;   // src/zipi8.vhd(327[13:15])
    
    wire ram_s_35_7, ram_s_32_3, ram_s_32_2, ram_s_32_1, ram_s_12_3, 
        ram_s_12_2, ram_s_36_2, ram_s_36_1, ram_s_37_4, ram_s_37_3, 
        ram_s_37_2, ram_s_39_5, ram_s_39_4, ram_s_39_3, ram_s_37_1, 
        ram_s_36_7, ram_s_37_0, ram_s_36_0, ram_s_6_4, ram_s_6_3, 
        ram_s_6_2, ram_s_6_1, ram_s_6_0, ram_s_5_7, ram_s_5_6, ram_s_5_5, 
        ram_s_5_4, ram_s_5_3, ram_s_5_2, ram_s_5_1, ram_s_5_0, ram_s_4_7, 
        ram_s_4_6, ram_s_4_5, ram_s_4_4, ram_s_4_3, ram_s_4_2, ram_s_4_1, 
        ram_s_4_0, ram_s_3_7, ram_s_3_6, ram_s_3_5, ram_s_35_6;
    wire [11:0]pc_value;   // src/program_counter.vhd(48[12:20])
    
    wire n893, ram_s_8_0, ram_s_13_7, ram_s_13_6, ram_s_13_5, ram_s_13_4, 
        ram_s_13_3, ram_s_13_2, ram_s_14_5, ram_s_14_4, ram_s_14_3, 
        ram_s_14_2, ram_s_14_1, ram_s_14_0, ram_s_14_7, ram_s_14_6, 
        ram_s_12_6, ram_s_13_1, ram_s_8_1, ram_s_13_0, ram_s_12_7, 
        ram_s_35_5, ram_s_12_5, ram_s_12_4, ram_s_12_1, ram_s_12_0, 
        ram_s_11_7, ram_s_11_6, ram_s_11_5, ram_s_11_4, ram_s_11_3, 
        ram_s_11_2, ram_s_11_1, ram_s_11_0, ram_s_3_4, ram_s_3_3, 
        ram_s_3_2, ram_s_3_1, ram_s_3_0, ram_s_2_7, ram_s_2_6, ram_s_2_5, 
        ram_s_2_4, ram_s_2_3, ram_s_2_2, ram_s_2_1, ram_s_2_0, ram_s_1_7, 
        ram_s_1_6, ram_s_1_5, ram_s_1_4, ram_s_1_3, ram_s_39_2, ram_s_39_1, 
        ram_s_39_0, ram_s_38_7, ram_s_38_6, ram_s_38_5, ram_s_38_4, 
        ram_s_38_3, ram_s_38_2, ram_s_38_1, ram_s_38_0, ram_s_37_7, 
        ram_s_37_6, ram_s_37_5, ram_s_40_7, ram_s_40_6, ram_s_35_4, 
        ram_s_40_5, ram_s_35_3, ram_s_35_0, ram_s_1_2, ram_s_1_1, 
        ram_s_1_0, ram_s_0_7, ram_s_0_5, ram_s_0_4, ram_s_0_3, ram_s_0_2, 
        ram_s_0_1, ram_s_0_0, ram_s_35_2, ram_s_40_4, ram_s_40_3, 
        ram_s_40_2, ram_s_35_1, ram_s_0_6, ram_s_40_1, ram_s_34_7, 
        ram_s_40_0, ram_s_34_6, ram_s_34_5, ram_s_34_4, ram_s_32_7, 
        ram_s_33_5, ram_s_7_7, ram_s_7_6, ram_s_34_1, ram_s_8_2, ram_s_34_0, 
        ram_s_33_7, ram_s_33_6, ram_s_34_3, ram_s_33_4, ram_s_33_3, 
        ram_s_33_2, ram_s_33_1, ram_s_33_0, ram_s_32_5, ram_s_32_4, 
        ram_s_7_5, ram_s_7_4, ram_s_7_3, ram_s_7_2, ram_s_7_1, ram_s_7_0, 
        ram_s_6_7, ram_s_6_6, ram_s_6_5, ram_s_34_2, ram_s_8_7, ram_s_8_6, 
        ram_s_8_5, ram_s_8_4, ram_s_8_3, ram_s_39_7, VCC_net, ram_s_39_6, 
        ram_s_44_2, ram_s_44_3, ram_s_44_4, ram_s_44_5, ram_s_44_6, 
        ram_s_44_7, ram_s_45_0, ram_s_45_1, ram_s_45_2, ram_s_45_3, 
        ram_s_45_4, ram_s_45_5, ram_s_45_6, ram_s_45_7, ram_s_47_0, 
        ram_s_47_1, ram_s_47_2, ram_s_47_3, ram_s_47_4, ram_s_47_5, 
        ram_s_47_6, ram_s_47_7, ram_s_57_0, ram_s_57_1, ram_s_57_2, 
        ram_s_57_3, ram_s_57_4, ram_s_57_5, ram_s_57_6, ram_s_57_7, 
        ram_s_58_0, ram_s_58_1, ram_s_58_2, ram_s_58_3, ram_s_58_4, 
        ram_s_58_5, ram_s_58_6, ram_s_58_7, ram_s_62_0, ram_s_62_1, 
        ram_s_62_2, ram_s_62_3, ram_s_62_4, ram_s_62_5, ram_s_62_6, 
        ram_s_62_7, ram_s_63_0, ram_s_63_1, ram_s_63_2, ram_s_63_3, 
        ram_s_63_4, ram_s_63_5, ram_s_63_6, ram_s_63_7, ram_s_64_0, 
        ram_s_64_1, ram_s_64_2, ram_s_64_3, ram_s_64_4, ram_s_64_5, 
        ram_s_64_6, ram_s_64_7, ram_s_65_0, ram_s_65_1, ram_s_65_2, 
        ram_s_65_3, ram_s_65_4, ram_s_65_5, ram_s_65_6, ram_s_65_7, 
        ram_s_66_0, ram_s_66_1, ram_s_66_2, ram_s_66_3, ram_s_66_4, 
        ram_s_66_5, ram_s_66_6, ram_s_66_7, ram_s_67_0, ram_s_67_1, 
        ram_s_67_2, ram_s_67_3, ram_s_67_4, ram_s_67_5, ram_s_67_6, 
        ram_s_67_7, ram_s_68_0, ram_s_68_1, ram_s_68_2, ram_s_68_3, 
        ram_s_68_4, ram_s_68_5, ram_s_68_6, ram_s_68_7, ram_s_69_0, 
        ram_s_69_1, ram_s_69_2, ram_s_69_3, ram_s_69_4, ram_s_69_5, 
        ram_s_69_6, ram_s_69_7, ram_s_70_0, ram_s_70_1, ram_s_70_2, 
        ram_s_70_3, ram_s_70_4, ram_s_70_5, ram_s_70_6, ram_s_70_7, 
        ram_s_71_0, ram_s_71_1, ram_s_71_2, ram_s_71_3, ram_s_71_4, 
        ram_s_71_5, ram_s_71_6, ram_s_71_7, ram_s_72_0, ram_s_72_1, 
        ram_s_72_2, ram_s_72_3, ram_s_72_4, ram_s_72_5, ram_s_72_6, 
        ram_s_72_7, ram_s_73_0, ram_s_73_1, ram_s_73_2, ram_s_73_3, 
        ram_s_73_4, ram_s_73_5, ram_s_73_6, ram_s_73_7, ram_s_74_0, 
        ram_s_74_1, ram_s_74_2, ram_s_74_3, ram_s_74_4, ram_s_74_5, 
        ram_s_74_6, ram_s_74_7, ram_s_75_0, ram_s_75_1, ram_s_75_2, 
        ram_s_75_3, ram_s_75_4, ram_s_75_5, ram_s_75_6, ram_s_75_7, 
        ram_s_81_0, ram_s_81_1, ram_s_81_2, ram_s_81_3, ram_s_81_4, 
        ram_s_81_5, ram_s_81_6, ram_s_81_7, ram_s_128_0, ram_s_128_1, 
        ram_s_128_2, ram_s_128_3, ram_s_128_4, ram_s_128_5, ram_s_128_6, 
        ram_s_128_7, ram_s_129_0, ram_s_129_1, ram_s_129_2, ram_s_129_3, 
        ram_s_129_4, ram_s_129_5, ram_s_129_6, ram_s_129_7, ram_s_130_0, 
        ram_s_130_1, ram_s_130_2, ram_s_130_3, ram_s_130_4, ram_s_130_5, 
        ram_s_130_6, ram_s_130_7, ram_s_131_0, ram_s_131_1, ram_s_131_2, 
        ram_s_131_3, ram_s_131_4, ram_s_131_5, ram_s_131_6, ram_s_131_7, 
        ram_s_132_0, ram_s_132_1, ram_s_132_2, ram_s_132_3, ram_s_132_4, 
        ram_s_132_5, ram_s_132_6, ram_s_132_7, ram_s_133_0, ram_s_133_1, 
        ram_s_133_2, ram_s_133_3, ram_s_133_4, ram_s_133_5, ram_s_133_6, 
        ram_s_133_7, ram_s_134_0, ram_s_134_1, ram_s_134_2, ram_s_134_3, 
        ram_s_134_4, ram_s_134_5, ram_s_134_6, ram_s_134_7, ram_s_135_0, 
        ram_s_135_1, ram_s_135_2, ram_s_135_3, ram_s_135_4, ram_s_135_5, 
        ram_s_135_6, ram_s_135_7, ram_s_136_0, ram_s_136_1, ram_s_136_2, 
        ram_s_136_3, ram_s_136_4, ram_s_136_5, ram_s_136_6, ram_s_136_7, 
        ram_s_139_0, ram_s_139_1, ram_s_139_2, ram_s_139_3, ram_s_139_4, 
        ram_s_139_5, ram_s_139_6, ram_s_139_7, ram_s_140_0, ram_s_140_1, 
        ram_s_140_2, ram_s_140_3, ram_s_140_4, ram_s_140_5, ram_s_140_6, 
        ram_s_140_7, ram_s_141_0, ram_s_141_1, ram_s_141_2, ram_s_141_3, 
        ram_s_141_4, ram_s_141_5, ram_s_141_6, ram_s_141_7, ram_s_142_0, 
        ram_s_142_1, ram_s_142_2, ram_s_142_3, ram_s_142_4, ram_s_142_5, 
        ram_s_142_6, ram_s_142_7, ram_s_160_0, ram_s_160_1, ram_s_160_2, 
        ram_s_160_3, ram_s_160_4, ram_s_160_5, ram_s_160_6, ram_s_160_7, 
        ram_s_161_0, ram_s_161_1, ram_s_161_2, ram_s_161_3, ram_s_161_4, 
        ram_s_161_5, ram_s_161_6, ram_s_161_7, ram_s_162_0, ram_s_162_1, 
        ram_s_162_2, ram_s_162_3, ram_s_162_4, ram_s_162_5, ram_s_162_6, 
        ram_s_162_7, ram_s_163_0, ram_s_163_1, ram_s_163_2, ram_s_163_3, 
        ram_s_163_4, ram_s_163_5, ram_s_163_6, ram_s_163_7, ram_s_164_0, 
        ram_s_164_1, ram_s_164_2, ram_s_164_3, ram_s_164_4, ram_s_164_5, 
        ram_s_164_6, ram_s_164_7, ram_s_165_0, ram_s_165_1, ram_s_165_2, 
        ram_s_165_3, ram_s_165_4, ram_s_165_5, ram_s_165_6, ram_s_165_7, 
        ram_s_166_0, ram_s_166_1, ram_s_166_2, ram_s_166_3, ram_s_166_4, 
        ram_s_166_5, ram_s_166_6, ram_s_166_7, ram_s_167_0, ram_s_167_1, 
        ram_s_167_2, ram_s_167_3, ram_s_167_4, ram_s_167_5, ram_s_167_6, 
        ram_s_167_7, ram_s_168_0, ram_s_168_1, ram_s_168_2, ram_s_168_3, 
        ram_s_168_4, ram_s_168_5, ram_s_168_6, ram_s_168_7, ram_s_171_0, 
        ram_s_171_1, ram_s_171_2, ram_s_171_3, ram_s_171_4, ram_s_171_5, 
        ram_s_171_6, ram_s_171_7, ram_s_172_0, ram_s_172_1, ram_s_172_2, 
        ram_s_172_3, ram_s_172_4, ram_s_172_5, ram_s_172_6, ram_s_172_7, 
        ram_s_173_0, ram_s_173_1, ram_s_173_2, ram_s_173_3, ram_s_173_4, 
        ram_s_173_5, ram_s_173_6, ram_s_173_7, ram_s_175_0, ram_s_175_1, 
        ram_s_175_2, ram_s_175_3, ram_s_175_4, ram_s_175_5, ram_s_175_6, 
        ram_s_175_7, ram_s_185_0, ram_s_185_1, ram_s_185_2, ram_s_185_3, 
        ram_s_185_4, ram_s_185_5, ram_s_185_6, ram_s_185_7, ram_s_186_0, 
        ram_s_186_1, ram_s_186_2, ram_s_186_3, ram_s_186_4, ram_s_186_5, 
        ram_s_186_6, ram_s_186_7, ram_s_190_0, ram_s_190_1, ram_s_190_2, 
        ram_s_190_3, ram_s_190_4, ram_s_190_5, ram_s_190_6, ram_s_190_7, 
        ram_s_191_0, ram_s_191_1, ram_s_191_2, ram_s_191_3, ram_s_191_4, 
        ram_s_191_5, ram_s_191_6, ram_s_191_7, ram_s_192_0, ram_s_192_1, 
        ram_s_192_2, ram_s_192_3, ram_s_192_4, ram_s_192_5, ram_s_192_6, 
        ram_s_192_7, ram_s_193_0, ram_s_193_1, ram_s_193_2, ram_s_193_3, 
        ram_s_193_4, ram_s_193_5, ram_s_193_6, ram_s_193_7, ram_s_194_0, 
        ram_s_194_1, ram_s_194_2, ram_s_194_3, ram_s_194_4, ram_s_194_5, 
        ram_s_194_6, ram_s_194_7, ram_s_195_0, ram_s_195_1, ram_s_195_2, 
        ram_s_195_3, ram_s_195_4, ram_s_195_5, ram_s_195_6, ram_s_195_7, 
        ram_s_196_0, ram_s_196_1, ram_s_196_2, ram_s_196_3, ram_s_196_4, 
        ram_s_196_5, ram_s_196_6, ram_s_196_7, ram_s_197_0, ram_s_197_1, 
        ram_s_197_2, ram_s_197_3, ram_s_197_4, ram_s_197_5, ram_s_197_6, 
        ram_s_197_7, ram_s_198_0, ram_s_198_1, ram_s_198_2, ram_s_198_3, 
        ram_s_198_4, ram_s_198_5, ram_s_198_6, ram_s_198_7, ram_s_199_0, 
        ram_s_199_1, ram_s_199_2, ram_s_199_3, ram_s_199_4, ram_s_199_5, 
        ram_s_199_6, ram_s_199_7, ram_s_200_0, ram_s_200_1, ram_s_200_2, 
        ram_s_200_3, ram_s_200_4, ram_s_200_5, ram_s_200_6, ram_s_200_7, 
        ram_s_201_0, ram_s_201_1, ram_s_201_2, ram_s_201_3, ram_s_201_4, 
        ram_s_201_5, ram_s_201_6, ram_s_201_7, ram_s_202_0, ram_s_202_1, 
        ram_s_202_2, ram_s_202_3, ram_s_202_4, ram_s_202_5, ram_s_202_6, 
        ram_s_202_7, ram_s_203_0, ram_s_203_1, ram_s_203_2, ram_s_203_3, 
        ram_s_203_4, ram_s_203_5, ram_s_203_6, ram_s_203_7, ram_s_209_0, 
        ram_s_209_1, ram_s_209_2, ram_s_209_3, ram_s_209_4, ram_s_209_5, 
        ram_s_209_6, ram_s_209_7, n48, n54, n55, n56, n57, n58, 
        n59, n60, n61, n62, n63, n64, n65, n66, n67, n71, 
        n72, n82, n84, n85, n86, n89, n90, n91, n92, n93, 
        n94, n95, n96, n97, n115, n116, n117, n118, n121, 
        n122, n123, n124, n125, n126, n127, n128, n129, n176, 
        n182, n183, n184, n185, n186, n187, n188, n189, n190, 
        n191, n192, n193, n194, n195, n199, n200, n210, n212, 
        n213, n214, n217, n218, n219, n220, n221, n222, n223, 
        n224, n225, n243, n244, n245, n246, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n2567, n2566, n2565, 
        n2564, n2563, n2562, n2561, n2560, n2519, n2518, n2517, 
        n2516, n2515, n2514, n2513, n2512, n2511, n2510, n2509, 
        n2508, n2507, n2506, n2505, n2504, n2503, n2502, n2501, 
        n2500, n2499, n2498, n2497, n2496, n2495, n2494, n2493, 
        n2492, n2491, n2490, n2489, n2488, n2487, n2486, n2485, 
        n2484, n2483, n2482, n2481, n2480, n2479, n2478, n2477, 
        n2476, n2475, n2474, n2473, n2472, n2471, n2470, n2469, 
        n2468, n2467, n2466, n2465, n2464, n2463, n2462, n2461, 
        n2460, n2459, n2458, n2457, n2456, n2455, n2454, n2453, 
        n2452, n2451, n2450, n2449, n2448, n2447, n2446, n2445, 
        n2444, n2443, n2442, n2441, n2440, n2439, n2438, n2437, 
        n2436, n2435, n2434, n2433, n2432, n2431, n2430, n2429, 
        n2428, n2427, n2426, n2425, n2424, n2423, n2422, n2421, 
        n2420, n2419, n2418, n2417, n2416, n2415, n2414, n2413, 
        n2412, n2411, n2410, n2409, n2408, n2383, n2382, n2381, 
        n2380, n2379, n2378, n2377, n2376, n2375, n2374, n2373, 
        n2372, n2371, n2370, n2369, n2368, n2295, n2294, n2293, 
        n2292, n2291, n2290, n2289, n2288, n2279, n2278, n2277, 
        n2276, n2275, n2274, n2273, n2272, n2271, n2270, n2269, 
        n2268, n2267, n2266, n2265, n2264, n2263, n2262, n2261, 
        n2260, n2259, n2258, n2257, n2256, n2239, n2238, n2237, 
        n2236, n2235, n2234, n2233, n2232, n2231, n2230, n2229, 
        n2228, n2227, n2226, n2225, n2224, n2223, n2222, n2221, 
        n2220, n2219, n2218, n2217, n2216, n2215, n2214, n2213, 
        n2212, n2211, n2210, n2209, n2208, n2207, n2206, n2205, 
        n2204, n2203, n2202, n2201, n2200, n2199, n2198, n2197, 
        n2196, n2195, n2194, n2193, n2192, n2191, n2190, n2189, 
        n2188, n2187, n2186, n2185, n2184, n2183, n2182, n2181, 
        n2180, n2179, n2178, n2177, n2176, n2175, n2174, n2173, 
        n2172, n2171, n2170, n2169, n2168, n2031, n2030, n2029, 
        n2028, n2027, n2026, n2025, n2024, n2023, n2022, n2021, 
        n2020, n2019, n2018, n2017, n2016, n2015, n2014, n2013, 
        n2012, n2011, n2010, n2009, n2008, n2007, n2006, n2005, 
        n2004, n2003, n2002, n2001, n2000, n1983, n1982, n1981, 
        n1980, n1979, n1978, n1977, n1976, n1975, n1974, n1973, 
        n1972, n1971, n1970, n1969, n1968, n1967, n1966, n1965, 
        n1964, n1963, n1962, n1961, n1960, n1959, n1958, n1957, 
        n1956, n1955, n1954, n1953, n1952, n1951, n1950, n1949, 
        n1948, n1947, n1946, n1945, n1944, n1943, n1942, n1941, 
        n1940, n1939, n1938, n1937, n1936, n1935, n1934, n1933, 
        n1932, n1931, n1930, n1929, n1928, n1927, n1926, n1925, 
        n1924, n1923, n1922, n1921, n1920, n1919, n1918, n1917, 
        n1916, n1915, n1914, n1913, n1912, n1543, n1542, n1541, 
        n1540, n1539, n1538, n1537, n1536, n1495, n1494, n1493, 
        n1492, n1491, n1490, n1489, n1488, n1487, n1486, n1485, 
        n1484, n1483, n1482, n1481, n1480, n1479, n1478, n1477, 
        n1476, n1475, n1474, n1473, n1472, n1471, n1470, n1469, 
        n1468, n1467, n1466, n1465, n1464, n1463, n1462, n1461, 
        n1460, n1459, n1458, n1457, n1456, n1455, n1454, n1453, 
        n1452, n1451, n1450, n1449, n1448, n1447, n1446, n1445, 
        n1444, n1443, n1442, n1441, n1440, n1439, n1438, n1437, 
        n1436, n1435, n1434, n1433, n1432, n1431, n1430, n1429, 
        n1428, n1427, n1426, n1425, n1424, n1423, n1422, n1421, 
        n1420, n1419, n1418, n1417, n1416, n1415, n1414, n1413, 
        n1412, n1411, n1410, n1409, n1408, n1407, n1406, n1405, 
        n1404, n1403, n1402, n1401, n1400, n1399, n1398, n1397, 
        n1396, n1395, n1394, n1393, n1392, n1391, n1390, n1389, 
        n1388, n1387, n1386, n1385, n1384, n1359, n1358, n1357, 
        n1356, n1355, n1354, n1353, n1352, n1351, n1350, n1349, 
        n1348, n1347, n1346, n1345, n1344, n1271, n1270, n1269, 
        n1268, n1267, n1266, n1265, n1264, n1255, n1254, n1253, 
        n1252, n1251, n1250, n1249, n1248, n1247, n1246, n1245, 
        n1244, n1243, n1242, n1241, n1240, n1239, n1238, n1237, 
        n1236, n1235, n1234, n1233, n1232, n1215, n1214, n1213, 
        n1212, n1211, n1210, n1209, n1208, n1207, n1206, n1205, 
        n1204, n1203, n1202, n1201, n1200, n1199, n1198, n1197, 
        n1196, n1195, n1194, n1193, n1192, n1191, n1190, n1189, 
        n1188, n1187, n1186, n1185, n1184, n1183, n1182, n1181, 
        n1180, n1179, n1178, n1177, n1176, n1175, n1174, n1173, 
        n1172, n1171, n1170, n1169, n1168, n1167, n1166, n1165, 
        n1164, n1163, n1162, n1161, n1160, n1159, n1158, n1157, 
        n1156, n1155, n1154, n1153, n1152, n1151, n1150, n1149, 
        n1148, n1147, n1146, n1145, n1144, n1051, n1047, n1046, 
        n1045, n1044, n1043, n1042, n1041, n1040, n1038, n1037, 
        n1036, n1035, n1034, n1033, n1032, n1031, n1030, n1029, 
        n1017, n1016, n1015, n1014, n1013, n1012, n1011, n1010, 
        n1009, n1008, n1007, n1006, n1005, n1004, n1003, n1002, 
        n1001, n998, n997, n996, n995, n994, n993, n992, n989, 
        n988, n987, n986, n985, n984, n983, n980, n979, n978, 
        n977, n976, n975, n974, n973, n972, n971, n970, n969, 
        n968, n967, n966, n965, n964, n963, n962, n961, n960, 
        n959, n958, n957, n952, n950, n946, n944, n941, n940, 
        n939, n938, n935, n934, n933, n932, n931, n930, n927, 
        n926, n925, n924, n923, n918, n917, n916, n8580, n765, 
        n911, n909, n908, n907, n906, n904, n901;
    
    VCC i2 (.Y(VCC_net));
    zipi8 processor_zipi8 (.CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .instruction({instruction}), 
          .wea({GND_net}), .\sx[7] (sx[7]), .\sx[6] (sx[6]), .\sx[5] (sx[5]), 
          .\sx[4] (sx[4]), .\register_vector[11] (register_vector[11]), 
          .\register_vector[10] (register_vector[10]), .\register_vector[9] (register_vector[9]), 
          .\register_vector[8] (register_vector[8]), .n8580(n8580), .bram_enable(bram_enable), 
          .\t_state[1] (t_state[1]), .internal_reset(internal_reset), .BTN1_c(BTN1_c), 
          .special_bit(special_bit), .address({Open_0, address[10:0]}), 
          .VCC_net(VCC_net), .ram_s_70_3(ram_s_70_3), .ram_s_71_3(ram_s_71_3), 
          .ram_s_69_3(ram_s_69_3), .ram_s_68_3(ram_s_68_3), .ram_s_34_7(ram_s_34_7), 
          .ram_s_35_7(ram_s_35_7), .ram_s_33_7(ram_s_33_7), .ram_s_32_7(ram_s_32_7), 
          .ram_s_11_6(ram_s_11_6), .ram_s_8_6(ram_s_8_6), .ram_s_62_4(ram_s_62_4), 
          .ram_s_63_4(ram_s_63_4), .ram_s_2_7(ram_s_2_7), .ram_s_3_7(ram_s_3_7), 
          .ram_s_1_7(ram_s_1_7), .ram_s_0_7(ram_s_0_7), .ram_s_66_4(ram_s_66_4), 
          .ram_s_67_4(ram_s_67_4), .ram_s_65_4(ram_s_65_4), .ram_s_64_4(ram_s_64_4), 
          .ram_s_142_3(ram_s_142_3), .ram_s_141_3(ram_s_141_3), .ram_s_140_3(ram_s_140_3), 
          .ram_s_209_3(ram_s_209_3), .ram_s_130_0(ram_s_130_0), .ram_s_131_0(ram_s_131_0), 
          .ram_s_129_0(ram_s_129_0), .ram_s_128_0(ram_s_128_0), .ram_s_70_4(ram_s_70_4), 
          .ram_s_71_4(ram_s_71_4), .ram_s_69_4(ram_s_69_4), .ram_s_68_4(ram_s_68_4), 
          .ram_s_171_5(ram_s_171_5), .ram_s_168_5(ram_s_168_5), .ram_s_14_6(ram_s_14_6), 
          .ram_s_13_6(ram_s_13_6), .ram_s_12_6(ram_s_12_6), .ram_s_202_1(ram_s_202_1), 
          .ram_s_203_1(ram_s_203_1), .ram_s_6_5(ram_s_6_5), .ram_s_7_5(ram_s_7_5), 
          .ram_s_14_5(ram_s_14_5), .ram_s_5_5(ram_s_5_5), .ram_s_4_5(ram_s_4_5), 
          .ram_s_13_5(ram_s_13_5), .ram_s_12_5(ram_s_12_5), .ram_s_43_2(ram_s_43_2), 
          .ram_s_2_0(ram_s_2_0), .ram_s_3_0(ram_s_3_0), .ram_s_2_1(ram_s_2_1), 
          .ram_s_3_1(ram_s_3_1), .ram_s_1_0(ram_s_1_0), .ram_s_0_0(ram_s_0_0), 
          .ram_s_66_0(ram_s_66_0), .ram_s_67_0(ram_s_67_0), .ram_s_34_1(ram_s_34_1), 
          .ram_s_35_1(ram_s_35_1), .ram_s_33_1(ram_s_33_1), .ram_s_32_1(ram_s_32_1), 
          .ram_s_201_1(ram_s_201_1), .ram_s_200_1(ram_s_200_1), .ram_s_1_1(ram_s_1_1), 
          .ram_s_0_1(ram_s_0_1), .ram_s_65_0(ram_s_65_0), .ram_s_64_0(ram_s_64_0), 
          .ram_s_11_2(ram_s_11_2), .ram_s_8_2(ram_s_8_2), .ram_s_38_0(ram_s_38_0), 
          .ram_s_39_0(ram_s_39_0), .ram_s_40_2(ram_s_40_2), .ram_s_74_7(ram_s_74_7), 
          .ram_s_75_7(ram_s_75_7), .ram_s_73_7(ram_s_73_7), .ram_s_72_7(ram_s_72_7), 
          .ram_s_130_7(ram_s_130_7), .ram_s_131_7(ram_s_131_7), .ram_s_129_7(ram_s_129_7), 
          .ram_s_128_7(ram_s_128_7), .ram_s_37_0(ram_s_37_0), .ram_s_36_0(ram_s_36_0), 
          .ram_s_142_5(ram_s_142_5), .ram_s_141_5(ram_s_141_5), .ram_s_140_5(ram_s_140_5), 
          .ram_s_62_0(ram_s_62_0), .ram_s_63_0(ram_s_63_0), .ram_s_194_1(ram_s_194_1), 
          .ram_s_195_1(ram_s_195_1), .ram_s_193_1(ram_s_193_1), .ram_s_192_1(ram_s_192_1), 
          .ram_s_74_4(ram_s_74_4), .ram_s_75_4(ram_s_75_4), .ram_s_73_4(ram_s_73_4), 
          .ram_s_72_4(ram_s_72_4), .ram_s_43_7(ram_s_43_7), .ram_s_40_7(ram_s_40_7), 
          .ram_s_74_2(ram_s_74_2), .ram_s_75_2(ram_s_75_2), .ram_s_73_2(ram_s_73_2), 
          .ram_s_72_2(ram_s_72_2), .ram_s_186_3(ram_s_186_3), .ram_s_185_3(ram_s_185_3), 
          .ram_s_190_2(ram_s_190_2), .ram_s_191_2(ram_s_191_2), .ram_s_43_1(ram_s_43_1), 
          .ram_s_40_1(ram_s_40_1), .ram_s_6_7(ram_s_6_7), .ram_s_7_7(ram_s_7_7), 
          .ram_s_134_0(ram_s_134_0), .ram_s_135_0(ram_s_135_0), .ram_s_5_7(ram_s_5_7), 
          .ram_s_4_7(ram_s_4_7), .ram_s_133_0(ram_s_133_0), .ram_s_132_0(ram_s_132_0), 
          .ram_s_34_2(ram_s_34_2), .ram_s_35_2(ram_s_35_2), .ram_s_58_5(ram_s_58_5), 
          .ram_s_58_0(ram_s_58_0), .ram_s_57_0(ram_s_57_0), .ram_s_139_0(ram_s_139_0), 
          .ram_s_136_0(ram_s_136_0), .ram_s_190_5(ram_s_190_5), .ram_s_191_5(ram_s_191_5), 
          .ram_s_57_5(ram_s_57_5), .ram_s_33_2(ram_s_33_2), .ram_s_32_2(ram_s_32_2), 
          .ram_s_142_7(ram_s_142_7), .ram_s_141_7(ram_s_141_7), .ram_s_140_7(ram_s_140_7), 
          .ram_s_81_5(ram_s_81_5), .ram_s_190_1(ram_s_190_1), .ram_s_191_1(ram_s_191_1), 
          .ram_s_139_1(ram_s_139_1), .ram_s_136_1(ram_s_136_1), .ram_s_38_7(ram_s_38_7), 
          .ram_s_39_7(ram_s_39_7), .ram_s_37_7(ram_s_37_7), .ram_s_36_7(ram_s_36_7), 
          .n893(n893), .ram_s_14_4(ram_s_14_4), .ram_s_190_7(ram_s_190_7), 
          .ram_s_191_7(ram_s_191_7), .ram_s_47_2(ram_s_47_2), .ram_s_45_2(ram_s_45_2), 
          .ram_s_44_2(ram_s_44_2), .ram_s_134_5(ram_s_134_5), .ram_s_135_5(ram_s_135_5), 
          .ram_s_133_5(ram_s_133_5), .ram_s_132_5(ram_s_132_5), .n2567(n2567), 
          .ram_s_209_7(ram_s_209_7), .n2566(n2566), .ram_s_209_6(ram_s_209_6), 
          .n2565(n2565), .ram_s_209_5(ram_s_209_5), .n2564(n2564), .ram_s_209_4(ram_s_209_4), 
          .n2563(n2563), .n2562(n2562), .ram_s_209_2(ram_s_209_2), .n2561(n2561), 
          .ram_s_209_1(ram_s_209_1), .n2560(n2560), .ram_s_209_0(ram_s_209_0), 
          .n2519(n2519), .ram_s_203_7(ram_s_203_7), .n2518(n2518), .ram_s_203_6(ram_s_203_6), 
          .n2517(n2517), .ram_s_203_5(ram_s_203_5), .n2516(n2516), .ram_s_203_4(ram_s_203_4), 
          .n2515(n2515), .ram_s_203_3(ram_s_203_3), .n2514(n2514), .ram_s_203_2(ram_s_203_2), 
          .n2513(n2513), .n2512(n2512), .ram_s_203_0(ram_s_203_0), .n2511(n2511), 
          .ram_s_202_7(ram_s_202_7), .n2510(n2510), .ram_s_202_6(ram_s_202_6), 
          .n2509(n2509), .ram_s_202_5(ram_s_202_5), .n2508(n2508), .ram_s_202_4(ram_s_202_4), 
          .n2507(n2507), .ram_s_202_3(ram_s_202_3), .n2506(n2506), .ram_s_202_2(ram_s_202_2), 
          .n2505(n2505), .n2504(n2504), .ram_s_202_0(ram_s_202_0), .n2503(n2503), 
          .ram_s_201_7(ram_s_201_7), .n2502(n2502), .ram_s_201_6(ram_s_201_6), 
          .n2501(n2501), .ram_s_201_5(ram_s_201_5), .n2500(n2500), .ram_s_201_4(ram_s_201_4), 
          .n2499(n2499), .ram_s_201_3(ram_s_201_3), .n2498(n2498), .ram_s_201_2(ram_s_201_2), 
          .n2497(n2497), .n2496(n2496), .ram_s_201_0(ram_s_201_0), .n2495(n2495), 
          .ram_s_200_7(ram_s_200_7), .n2494(n2494), .ram_s_200_6(ram_s_200_6), 
          .n2493(n2493), .ram_s_200_5(ram_s_200_5), .n2492(n2492), .ram_s_200_4(ram_s_200_4), 
          .n2491(n2491), .ram_s_200_3(ram_s_200_3), .n2490(n2490), .ram_s_200_2(ram_s_200_2), 
          .n2489(n2489), .n2488(n2488), .ram_s_200_0(ram_s_200_0), .n2487(n2487), 
          .ram_s_199_7(ram_s_199_7), .n2486(n2486), .ram_s_199_6(ram_s_199_6), 
          .n2485(n2485), .ram_s_199_5(ram_s_199_5), .n2484(n2484), .ram_s_199_4(ram_s_199_4), 
          .n2483(n2483), .ram_s_199_3(ram_s_199_3), .n2482(n2482), .ram_s_199_2(ram_s_199_2), 
          .n2481(n2481), .ram_s_199_1(ram_s_199_1), .n2480(n2480), .ram_s_199_0(ram_s_199_0), 
          .n2479(n2479), .ram_s_198_7(ram_s_198_7), .n2478(n2478), .ram_s_198_6(ram_s_198_6), 
          .n2477(n2477), .ram_s_198_5(ram_s_198_5), .n2476(n2476), .ram_s_198_4(ram_s_198_4), 
          .n2475(n2475), .ram_s_198_3(ram_s_198_3), .n2474(n2474), .ram_s_198_2(ram_s_198_2), 
          .n2473(n2473), .ram_s_198_1(ram_s_198_1), .n2472(n2472), .ram_s_198_0(ram_s_198_0), 
          .n2471(n2471), .ram_s_197_7(ram_s_197_7), .n2470(n2470), .ram_s_197_6(ram_s_197_6), 
          .n2469(n2469), .ram_s_197_5(ram_s_197_5), .n2468(n2468), .ram_s_197_4(ram_s_197_4), 
          .n2467(n2467), .ram_s_197_3(ram_s_197_3), .n2466(n2466), .ram_s_197_2(ram_s_197_2), 
          .n2465(n2465), .ram_s_197_1(ram_s_197_1), .n2464(n2464), .ram_s_197_0(ram_s_197_0), 
          .n2463(n2463), .ram_s_196_7(ram_s_196_7), .n2462(n2462), .ram_s_196_6(ram_s_196_6), 
          .n2461(n2461), .ram_s_196_5(ram_s_196_5), .n2460(n2460), .ram_s_196_4(ram_s_196_4), 
          .n2459(n2459), .ram_s_196_3(ram_s_196_3), .n2458(n2458), .ram_s_196_2(ram_s_196_2), 
          .n2457(n2457), .ram_s_196_1(ram_s_196_1), .n2456(n2456), .ram_s_196_0(ram_s_196_0), 
          .n2455(n2455), .ram_s_195_7(ram_s_195_7), .n2454(n2454), .ram_s_195_6(ram_s_195_6), 
          .n2453(n2453), .ram_s_195_5(ram_s_195_5), .n2452(n2452), .ram_s_195_4(ram_s_195_4), 
          .n2451(n2451), .ram_s_195_3(ram_s_195_3), .n2450(n2450), .ram_s_195_2(ram_s_195_2), 
          .n2449(n2449), .n2448(n2448), .ram_s_195_0(ram_s_195_0), .n2447(n2447), 
          .ram_s_194_7(ram_s_194_7), .n2446(n2446), .ram_s_194_6(ram_s_194_6), 
          .n2445(n2445), .ram_s_194_5(ram_s_194_5), .n2444(n2444), .ram_s_194_4(ram_s_194_4), 
          .n2443(n2443), .ram_s_194_3(ram_s_194_3), .n2442(n2442), .ram_s_194_2(ram_s_194_2), 
          .n2441(n2441), .n2440(n2440), .ram_s_194_0(ram_s_194_0), .n2439(n2439), 
          .ram_s_193_7(ram_s_193_7), .n2438(n2438), .ram_s_193_6(ram_s_193_6), 
          .n2437(n2437), .ram_s_193_5(ram_s_193_5), .n2436(n2436), .ram_s_193_4(ram_s_193_4), 
          .n2435(n2435), .ram_s_193_3(ram_s_193_3), .n2434(n2434), .ram_s_193_2(ram_s_193_2), 
          .n2433(n2433), .n2432(n2432), .ram_s_193_0(ram_s_193_0), .n2431(n2431), 
          .ram_s_192_7(ram_s_192_7), .n2430(n2430), .ram_s_192_6(ram_s_192_6), 
          .n2429(n2429), .ram_s_192_5(ram_s_192_5), .n2428(n2428), .ram_s_192_4(ram_s_192_4), 
          .n2427(n2427), .ram_s_192_3(ram_s_192_3), .n2426(n2426), .ram_s_192_2(ram_s_192_2), 
          .n2425(n2425), .n2424(n2424), .ram_s_192_0(ram_s_192_0), .n2423(n2423), 
          .n2422(n2422), .ram_s_191_6(ram_s_191_6), .n2421(n2421), .n2420(n2420), 
          .ram_s_191_4(ram_s_191_4), .n2419(n2419), .ram_s_191_3(ram_s_191_3), 
          .n2418(n2418), .n2417(n2417), .n2416(n2416), .ram_s_191_0(ram_s_191_0), 
          .n2415(n2415), .n2414(n2414), .ram_s_190_6(ram_s_190_6), .n2413(n2413), 
          .n2412(n2412), .ram_s_190_4(ram_s_190_4), .n2411(n2411), .ram_s_190_3(ram_s_190_3), 
          .n2410(n2410), .n2409(n2409), .n2408(n2408), .ram_s_190_0(ram_s_190_0), 
          .n2383(n2383), .ram_s_186_7(ram_s_186_7), .n2382(n2382), .ram_s_186_6(ram_s_186_6), 
          .n2381(n2381), .ram_s_186_5(ram_s_186_5), .n2380(n2380), .ram_s_186_4(ram_s_186_4), 
          .n2379(n2379), .n2378(n2378), .ram_s_186_2(ram_s_186_2), .n2377(n2377), 
          .ram_s_186_1(ram_s_186_1), .n2376(n2376), .ram_s_186_0(ram_s_186_0), 
          .n2375(n2375), .ram_s_185_7(ram_s_185_7), .n2374(n2374), .ram_s_185_6(ram_s_185_6), 
          .n2373(n2373), .ram_s_185_5(ram_s_185_5), .n2372(n2372), .ram_s_185_4(ram_s_185_4), 
          .n2371(n2371), .n2370(n2370), .ram_s_185_2(ram_s_185_2), .n2369(n2369), 
          .ram_s_185_1(ram_s_185_1), .n2368(n2368), .ram_s_185_0(ram_s_185_0), 
          .n2295(n2295), .ram_s_175_7(ram_s_175_7), .n2294(n2294), .ram_s_175_6(ram_s_175_6), 
          .n2293(n2293), .ram_s_175_5(ram_s_175_5), .n2292(n2292), .ram_s_175_4(ram_s_175_4), 
          .n2291(n2291), .ram_s_175_3(ram_s_175_3), .n2290(n2290), .ram_s_175_2(ram_s_175_2), 
          .n2289(n2289), .ram_s_175_1(ram_s_175_1), .n2288(n2288), .ram_s_175_0(ram_s_175_0), 
          .n2279(n2279), .ram_s_173_7(ram_s_173_7), .n2278(n2278), .ram_s_173_6(ram_s_173_6), 
          .n2277(n2277), .ram_s_173_5(ram_s_173_5), .n2276(n2276), .ram_s_173_4(ram_s_173_4), 
          .n2275(n2275), .ram_s_173_3(ram_s_173_3), .n2274(n2274), .ram_s_173_2(ram_s_173_2), 
          .n2273(n2273), .ram_s_173_1(ram_s_173_1), .n2272(n2272), .ram_s_173_0(ram_s_173_0), 
          .n2271(n2271), .ram_s_172_7(ram_s_172_7), .n2270(n2270), .ram_s_172_6(ram_s_172_6), 
          .n2269(n2269), .ram_s_172_5(ram_s_172_5), .n2268(n2268), .ram_s_172_4(ram_s_172_4), 
          .n2267(n2267), .ram_s_172_3(ram_s_172_3), .n2266(n2266), .ram_s_172_2(ram_s_172_2), 
          .n2265(n2265), .ram_s_172_1(ram_s_172_1), .n2264(n2264), .ram_s_172_0(ram_s_172_0), 
          .n2263(n2263), .ram_s_171_7(ram_s_171_7), .n2262(n2262), .ram_s_171_6(ram_s_171_6), 
          .n2261(n2261), .n2260(n2260), .ram_s_171_4(ram_s_171_4), .n2259(n2259), 
          .ram_s_171_3(ram_s_171_3), .n2258(n2258), .ram_s_171_2(ram_s_171_2), 
          .n2257(n2257), .ram_s_171_1(ram_s_171_1), .n2256(n2256), .ram_s_171_0(ram_s_171_0), 
          .n2239(n2239), .ram_s_168_7(ram_s_168_7), .n2238(n2238), .ram_s_168_6(ram_s_168_6), 
          .n2237(n2237), .n2236(n2236), .ram_s_168_4(ram_s_168_4), .n2235(n2235), 
          .ram_s_168_3(ram_s_168_3), .n2234(n2234), .ram_s_168_2(ram_s_168_2), 
          .n2233(n2233), .ram_s_168_1(ram_s_168_1), .n2232(n2232), .ram_s_168_0(ram_s_168_0), 
          .n2231(n2231), .ram_s_167_7(ram_s_167_7), .n2230(n2230), .ram_s_167_6(ram_s_167_6), 
          .n2229(n2229), .ram_s_167_5(ram_s_167_5), .n2228(n2228), .ram_s_167_4(ram_s_167_4), 
          .n2227(n2227), .ram_s_167_3(ram_s_167_3), .n2226(n2226), .ram_s_167_2(ram_s_167_2), 
          .n2225(n2225), .ram_s_167_1(ram_s_167_1), .n2224(n2224), .ram_s_167_0(ram_s_167_0), 
          .n2223(n2223), .ram_s_166_7(ram_s_166_7), .n2222(n2222), .ram_s_166_6(ram_s_166_6), 
          .n2221(n2221), .ram_s_166_5(ram_s_166_5), .n2220(n2220), .ram_s_166_4(ram_s_166_4), 
          .n2219(n2219), .ram_s_166_3(ram_s_166_3), .n2218(n2218), .ram_s_166_2(ram_s_166_2), 
          .n2217(n2217), .ram_s_166_1(ram_s_166_1), .n2216(n2216), .ram_s_166_0(ram_s_166_0), 
          .n2215(n2215), .ram_s_165_7(ram_s_165_7), .n2214(n2214), .ram_s_165_6(ram_s_165_6), 
          .n2213(n2213), .ram_s_165_5(ram_s_165_5), .n2212(n2212), .ram_s_165_4(ram_s_165_4), 
          .n2211(n2211), .ram_s_165_3(ram_s_165_3), .n2210(n2210), .ram_s_165_2(ram_s_165_2), 
          .n2209(n2209), .ram_s_165_1(ram_s_165_1), .n2208(n2208), .ram_s_165_0(ram_s_165_0), 
          .n2207(n2207), .ram_s_164_7(ram_s_164_7), .n2206(n2206), .ram_s_164_6(ram_s_164_6), 
          .n2205(n2205), .ram_s_164_5(ram_s_164_5), .n2204(n2204), .ram_s_164_4(ram_s_164_4), 
          .n2203(n2203), .ram_s_164_3(ram_s_164_3), .n2202(n2202), .ram_s_164_2(ram_s_164_2), 
          .n2201(n2201), .ram_s_164_1(ram_s_164_1), .n2200(n2200), .ram_s_164_0(ram_s_164_0), 
          .n2199(n2199), .ram_s_163_7(ram_s_163_7), .n2198(n2198), .ram_s_163_6(ram_s_163_6), 
          .n2197(n2197), .ram_s_163_5(ram_s_163_5), .n2196(n2196), .ram_s_163_4(ram_s_163_4), 
          .n2195(n2195), .ram_s_163_3(ram_s_163_3), .n2194(n2194), .ram_s_163_2(ram_s_163_2), 
          .n2193(n2193), .ram_s_163_1(ram_s_163_1), .n2192(n2192), .ram_s_163_0(ram_s_163_0), 
          .n2191(n2191), .ram_s_162_7(ram_s_162_7), .n2190(n2190), .ram_s_162_6(ram_s_162_6), 
          .n2189(n2189), .ram_s_162_5(ram_s_162_5), .n2188(n2188), .ram_s_162_4(ram_s_162_4), 
          .n2187(n2187), .ram_s_162_3(ram_s_162_3), .n2186(n2186), .ram_s_162_2(ram_s_162_2), 
          .n2185(n2185), .ram_s_162_1(ram_s_162_1), .n2184(n2184), .ram_s_162_0(ram_s_162_0), 
          .n2183(n2183), .ram_s_161_7(ram_s_161_7), .n2182(n2182), .ram_s_161_6(ram_s_161_6), 
          .n2181(n2181), .ram_s_161_5(ram_s_161_5), .n2180(n2180), .ram_s_161_4(ram_s_161_4), 
          .n2179(n2179), .ram_s_161_3(ram_s_161_3), .n2178(n2178), .ram_s_161_2(ram_s_161_2), 
          .n2177(n2177), .ram_s_161_1(ram_s_161_1), .n2176(n2176), .ram_s_161_0(ram_s_161_0), 
          .n2175(n2175), .ram_s_160_7(ram_s_160_7), .n2174(n2174), .ram_s_160_6(ram_s_160_6), 
          .n2173(n2173), .ram_s_160_5(ram_s_160_5), .n2172(n2172), .ram_s_160_4(ram_s_160_4), 
          .n2171(n2171), .ram_s_160_3(ram_s_160_3), .n2170(n2170), .ram_s_160_2(ram_s_160_2), 
          .n2169(n2169), .ram_s_160_1(ram_s_160_1), .n2168(n2168), .ram_s_160_0(ram_s_160_0), 
          .n2031(n2031), .n2030(n2030), .ram_s_142_6(ram_s_142_6), .n2029(n2029), 
          .n2028(n2028), .ram_s_142_4(ram_s_142_4), .n2027(n2027), .n2026(n2026), 
          .ram_s_142_2(ram_s_142_2), .n2025(n2025), .ram_s_142_1(ram_s_142_1), 
          .n2024(n2024), .ram_s_142_0(ram_s_142_0), .n2023(n2023), .n2022(n2022), 
          .ram_s_141_6(ram_s_141_6), .n2021(n2021), .n2020(n2020), .ram_s_141_4(ram_s_141_4), 
          .n2019(n2019), .n2018(n2018), .ram_s_141_2(ram_s_141_2), .n2017(n2017), 
          .ram_s_141_1(ram_s_141_1), .n2016(n2016), .ram_s_141_0(ram_s_141_0), 
          .n2015(n2015), .n2014(n2014), .ram_s_140_6(ram_s_140_6), .n2013(n2013), 
          .n2012(n2012), .ram_s_140_4(ram_s_140_4), .n2011(n2011), .n2010(n2010), 
          .ram_s_140_2(ram_s_140_2), .n2009(n2009), .ram_s_140_1(ram_s_140_1), 
          .n2008(n2008), .ram_s_140_0(ram_s_140_0), .n2007(n2007), .ram_s_139_7(ram_s_139_7), 
          .n2006(n2006), .ram_s_139_6(ram_s_139_6), .n2005(n2005), .ram_s_139_5(ram_s_139_5), 
          .n2004(n2004), .ram_s_139_4(ram_s_139_4), .n2003(n2003), .ram_s_139_3(ram_s_139_3), 
          .n2002(n2002), .ram_s_139_2(ram_s_139_2), .n2001(n2001), .n2000(n2000), 
          .n1983(n1983), .ram_s_136_7(ram_s_136_7), .n1982(n1982), .ram_s_136_6(ram_s_136_6), 
          .n1981(n1981), .ram_s_136_5(ram_s_136_5), .n1980(n1980), .ram_s_136_4(ram_s_136_4), 
          .n1979(n1979), .ram_s_136_3(ram_s_136_3), .n1978(n1978), .ram_s_136_2(ram_s_136_2), 
          .n1977(n1977), .n1976(n1976), .n1975(n1975), .ram_s_135_7(ram_s_135_7), 
          .n1974(n1974), .ram_s_135_6(ram_s_135_6), .n1973(n1973), .n1972(n1972), 
          .ram_s_135_4(ram_s_135_4), .n1971(n1971), .ram_s_135_3(ram_s_135_3), 
          .n1970(n1970), .ram_s_135_2(ram_s_135_2), .n1969(n1969), .ram_s_135_1(ram_s_135_1), 
          .n1968(n1968), .n1967(n1967), .ram_s_134_7(ram_s_134_7), .n1966(n1966), 
          .ram_s_134_6(ram_s_134_6), .n1965(n1965), .n1964(n1964), .ram_s_134_4(ram_s_134_4), 
          .n1963(n1963), .ram_s_134_3(ram_s_134_3), .n1962(n1962), .ram_s_134_2(ram_s_134_2), 
          .n1961(n1961), .ram_s_134_1(ram_s_134_1), .n1960(n1960), .n1959(n1959), 
          .ram_s_133_7(ram_s_133_7), .n1958(n1958), .ram_s_133_6(ram_s_133_6), 
          .n1957(n1957), .n1956(n1956), .ram_s_133_4(ram_s_133_4), .n1955(n1955), 
          .ram_s_133_3(ram_s_133_3), .n1954(n1954), .ram_s_133_2(ram_s_133_2), 
          .n1953(n1953), .ram_s_133_1(ram_s_133_1), .n1952(n1952), .n1951(n1951), 
          .ram_s_132_7(ram_s_132_7), .n1950(n1950), .ram_s_132_6(ram_s_132_6), 
          .n1949(n1949), .n1948(n1948), .ram_s_132_4(ram_s_132_4), .n1947(n1947), 
          .ram_s_132_3(ram_s_132_3), .n1946(n1946), .ram_s_132_2(ram_s_132_2), 
          .n1945(n1945), .ram_s_132_1(ram_s_132_1), .n1944(n1944), .n1943(n1943), 
          .n1942(n1942), .ram_s_131_6(ram_s_131_6), .n1941(n1941), .ram_s_131_5(ram_s_131_5), 
          .n1940(n1940), .ram_s_131_4(ram_s_131_4), .n1939(n1939), .ram_s_131_3(ram_s_131_3), 
          .n1938(n1938), .ram_s_131_2(ram_s_131_2), .n1937(n1937), .ram_s_131_1(ram_s_131_1), 
          .n1936(n1936), .n1935(n1935), .n1934(n1934), .ram_s_130_6(ram_s_130_6), 
          .n1933(n1933), .ram_s_130_5(ram_s_130_5), .n1932(n1932), .ram_s_130_4(ram_s_130_4), 
          .n1931(n1931), .ram_s_130_3(ram_s_130_3), .n1930(n1930), .ram_s_130_2(ram_s_130_2), 
          .n1929(n1929), .ram_s_130_1(ram_s_130_1), .n1928(n1928), .n1927(n1927), 
          .n1926(n1926), .ram_s_129_6(ram_s_129_6), .n1925(n1925), .ram_s_129_5(ram_s_129_5), 
          .n1924(n1924), .ram_s_129_4(ram_s_129_4), .n1923(n1923), .ram_s_129_3(ram_s_129_3), 
          .n1922(n1922), .ram_s_129_2(ram_s_129_2), .n1921(n1921), .ram_s_129_1(ram_s_129_1), 
          .n1920(n1920), .n1919(n1919), .n1918(n1918), .ram_s_128_6(ram_s_128_6), 
          .n1917(n1917), .ram_s_128_5(ram_s_128_5), .n1916(n1916), .ram_s_128_4(ram_s_128_4), 
          .n1915(n1915), .ram_s_128_3(ram_s_128_3), .n1914(n1914), .ram_s_128_2(ram_s_128_2), 
          .n1913(n1913), .ram_s_128_1(ram_s_128_1), .n1912(n1912), .n1543(n1543), 
          .ram_s_81_7(ram_s_81_7), .n1542(n1542), .ram_s_81_6(ram_s_81_6), 
          .n1541(n1541), .n1540(n1540), .ram_s_81_4(ram_s_81_4), .n1539(n1539), 
          .ram_s_81_3(ram_s_81_3), .n1538(n1538), .ram_s_81_2(ram_s_81_2), 
          .n1537(n1537), .ram_s_81_1(ram_s_81_1), .n1536(n1536), .ram_s_81_0(ram_s_81_0), 
          .n1495(n1495), .n1494(n1494), .ram_s_75_6(ram_s_75_6), .n1493(n1493), 
          .ram_s_75_5(ram_s_75_5), .n1492(n1492), .n1491(n1491), .ram_s_75_3(ram_s_75_3), 
          .n1490(n1490), .n1489(n1489), .ram_s_75_1(ram_s_75_1), .n1488(n1488), 
          .ram_s_75_0(ram_s_75_0), .n1487(n1487), .n1486(n1486), .ram_s_74_6(ram_s_74_6), 
          .n1485(n1485), .ram_s_74_5(ram_s_74_5), .n1484(n1484), .n1483(n1483), 
          .ram_s_74_3(ram_s_74_3), .n1482(n1482), .n1481(n1481), .ram_s_74_1(ram_s_74_1), 
          .n1480(n1480), .ram_s_74_0(ram_s_74_0), .n1479(n1479), .n1478(n1478), 
          .ram_s_73_6(ram_s_73_6), .n1477(n1477), .ram_s_73_5(ram_s_73_5), 
          .n1476(n1476), .n1475(n1475), .ram_s_73_3(ram_s_73_3), .n1474(n1474), 
          .n1473(n1473), .ram_s_73_1(ram_s_73_1), .n1472(n1472), .ram_s_73_0(ram_s_73_0), 
          .n1471(n1471), .n1470(n1470), .ram_s_72_6(ram_s_72_6), .n1469(n1469), 
          .ram_s_72_5(ram_s_72_5), .n1468(n1468), .n1467(n1467), .ram_s_72_3(ram_s_72_3), 
          .n1466(n1466), .n1465(n1465), .ram_s_72_1(ram_s_72_1), .n1464(n1464), 
          .ram_s_72_0(ram_s_72_0), .n1463(n1463), .ram_s_71_7(ram_s_71_7), 
          .n1462(n1462), .ram_s_71_6(ram_s_71_6), .n1461(n1461), .ram_s_71_5(ram_s_71_5), 
          .n1460(n1460), .n1459(n1459), .n1458(n1458), .ram_s_71_2(ram_s_71_2), 
          .n1457(n1457), .ram_s_71_1(ram_s_71_1), .n1456(n1456), .ram_s_71_0(ram_s_71_0), 
          .n1455(n1455), .ram_s_70_7(ram_s_70_7), .n1454(n1454), .ram_s_70_6(ram_s_70_6), 
          .n1453(n1453), .ram_s_70_5(ram_s_70_5), .n1452(n1452), .n1451(n1451), 
          .n1450(n1450), .ram_s_70_2(ram_s_70_2), .n1449(n1449), .ram_s_70_1(ram_s_70_1), 
          .n1448(n1448), .ram_s_70_0(ram_s_70_0), .n1447(n1447), .ram_s_69_7(ram_s_69_7), 
          .n1446(n1446), .ram_s_69_6(ram_s_69_6), .n1445(n1445), .ram_s_69_5(ram_s_69_5), 
          .n1444(n1444), .n1443(n1443), .n1442(n1442), .ram_s_69_2(ram_s_69_2), 
          .n1441(n1441), .ram_s_69_1(ram_s_69_1), .n1440(n1440), .ram_s_69_0(ram_s_69_0), 
          .n1439(n1439), .ram_s_68_7(ram_s_68_7), .n1438(n1438), .ram_s_68_6(ram_s_68_6), 
          .n1437(n1437), .ram_s_68_5(ram_s_68_5), .n1436(n1436), .n1435(n1435), 
          .n1434(n1434), .ram_s_68_2(ram_s_68_2), .n1433(n1433), .ram_s_68_1(ram_s_68_1), 
          .n1432(n1432), .ram_s_68_0(ram_s_68_0), .n1431(n1431), .ram_s_67_7(ram_s_67_7), 
          .n1430(n1430), .ram_s_67_6(ram_s_67_6), .n1429(n1429), .ram_s_67_5(ram_s_67_5), 
          .n1428(n1428), .n1427(n1427), .ram_s_67_3(ram_s_67_3), .n1426(n1426), 
          .ram_s_67_2(ram_s_67_2), .n1425(n1425), .ram_s_67_1(ram_s_67_1), 
          .n1424(n1424), .n1423(n1423), .ram_s_66_7(ram_s_66_7), .n1422(n1422), 
          .ram_s_66_6(ram_s_66_6), .n1421(n1421), .ram_s_66_5(ram_s_66_5), 
          .n1420(n1420), .n1419(n1419), .ram_s_66_3(ram_s_66_3), .n1418(n1418), 
          .ram_s_66_2(ram_s_66_2), .n1417(n1417), .ram_s_66_1(ram_s_66_1), 
          .n1416(n1416), .n1415(n1415), .ram_s_65_7(ram_s_65_7), .n1414(n1414), 
          .ram_s_65_6(ram_s_65_6), .n1413(n1413), .ram_s_65_5(ram_s_65_5), 
          .n1412(n1412), .n1411(n1411), .ram_s_65_3(ram_s_65_3), .n1410(n1410), 
          .ram_s_65_2(ram_s_65_2), .n1409(n1409), .ram_s_65_1(ram_s_65_1), 
          .n1408(n1408), .n1407(n1407), .ram_s_64_7(ram_s_64_7), .n1406(n1406), 
          .ram_s_64_6(ram_s_64_6), .n1405(n1405), .ram_s_64_5(ram_s_64_5), 
          .n1404(n1404), .n1403(n1403), .ram_s_64_3(ram_s_64_3), .n1402(n1402), 
          .ram_s_64_2(ram_s_64_2), .n1401(n1401), .ram_s_64_1(ram_s_64_1), 
          .n1400(n1400), .n1399(n1399), .ram_s_63_7(ram_s_63_7), .n1398(n1398), 
          .ram_s_63_6(ram_s_63_6), .n1397(n1397), .ram_s_63_5(ram_s_63_5), 
          .n1396(n1396), .n1395(n1395), .ram_s_63_3(ram_s_63_3), .n1394(n1394), 
          .ram_s_63_2(ram_s_63_2), .n1393(n1393), .ram_s_63_1(ram_s_63_1), 
          .n1392(n1392), .n1391(n1391), .ram_s_62_7(ram_s_62_7), .n1390(n1390), 
          .ram_s_62_6(ram_s_62_6), .n1389(n1389), .ram_s_62_5(ram_s_62_5), 
          .n1388(n1388), .n1387(n1387), .ram_s_62_3(ram_s_62_3), .n1386(n1386), 
          .ram_s_62_2(ram_s_62_2), .n1385(n1385), .ram_s_62_1(ram_s_62_1), 
          .n1384(n1384), .n1359(n1359), .ram_s_58_7(ram_s_58_7), .n1358(n1358), 
          .ram_s_58_6(ram_s_58_6), .n1357(n1357), .n1356(n1356), .ram_s_58_4(ram_s_58_4), 
          .n1355(n1355), .ram_s_58_3(ram_s_58_3), .n1354(n1354), .ram_s_58_2(ram_s_58_2), 
          .n1353(n1353), .ram_s_58_1(ram_s_58_1), .n1352(n1352), .n1351(n1351), 
          .ram_s_57_7(ram_s_57_7), .n1350(n1350), .ram_s_57_6(ram_s_57_6), 
          .n1349(n1349), .n1348(n1348), .ram_s_57_4(ram_s_57_4), .n1347(n1347), 
          .ram_s_57_3(ram_s_57_3), .n1346(n1346), .ram_s_57_2(ram_s_57_2), 
          .n1345(n1345), .ram_s_57_1(ram_s_57_1), .n1344(n1344), .n1271(n1271), 
          .ram_s_47_7(ram_s_47_7), .n1270(n1270), .ram_s_47_6(ram_s_47_6), 
          .n1269(n1269), .ram_s_47_5(ram_s_47_5), .n1268(n1268), .ram_s_47_4(ram_s_47_4), 
          .n1267(n1267), .ram_s_47_3(ram_s_47_3), .n1266(n1266), .n1265(n1265), 
          .ram_s_47_1(ram_s_47_1), .n1264(n1264), .ram_s_47_0(ram_s_47_0), 
          .n1255(n1255), .ram_s_45_7(ram_s_45_7), .n1254(n1254), .ram_s_45_6(ram_s_45_6), 
          .n1253(n1253), .ram_s_45_5(ram_s_45_5), .n1252(n1252), .ram_s_45_4(ram_s_45_4), 
          .n1251(n1251), .ram_s_45_3(ram_s_45_3), .n1250(n1250), .n1249(n1249), 
          .ram_s_45_1(ram_s_45_1), .n1248(n1248), .ram_s_45_0(ram_s_45_0), 
          .n1247(n1247), .ram_s_44_7(ram_s_44_7), .n1246(n1246), .ram_s_44_6(ram_s_44_6), 
          .n1245(n1245), .ram_s_44_5(ram_s_44_5), .n1244(n1244), .ram_s_44_4(ram_s_44_4), 
          .n1243(n1243), .ram_s_44_3(ram_s_44_3), .n1242(n1242), .n1241(n1241), 
          .ram_s_44_1(ram_s_44_1), .n1240(n1240), .ram_s_44_0(ram_s_44_0), 
          .n1239(n1239), .n1238(n1238), .ram_s_43_6(ram_s_43_6), .n1237(n1237), 
          .ram_s_43_5(ram_s_43_5), .n1236(n1236), .ram_s_43_4(ram_s_43_4), 
          .n1235(n1235), .ram_s_43_3(ram_s_43_3), .n1234(n1234), .n1233(n1233), 
          .n1232(n1232), .ram_s_43_0(ram_s_43_0), .n1215(n1215), .n1214(n1214), 
          .ram_s_40_6(ram_s_40_6), .n1213(n1213), .ram_s_40_5(ram_s_40_5), 
          .n1212(n1212), .ram_s_40_4(ram_s_40_4), .n1211(n1211), .ram_s_40_3(ram_s_40_3), 
          .n1210(n1210), .n1209(n1209), .n1208(n1208), .ram_s_40_0(ram_s_40_0), 
          .n1207(n1207), .n1206(n1206), .ram_s_39_6(ram_s_39_6), .n1205(n1205), 
          .ram_s_39_5(ram_s_39_5), .n1204(n1204), .ram_s_39_4(ram_s_39_4), 
          .n1203(n1203), .ram_s_39_3(ram_s_39_3), .n1202(n1202), .ram_s_39_2(ram_s_39_2), 
          .n1201(n1201), .ram_s_39_1(ram_s_39_1), .n1200(n1200), .n1199(n1199), 
          .n1198(n1198), .ram_s_38_6(ram_s_38_6), .n1197(n1197), .ram_s_38_5(ram_s_38_5), 
          .n1196(n1196), .ram_s_38_4(ram_s_38_4), .n1195(n1195), .ram_s_38_3(ram_s_38_3), 
          .n1194(n1194), .ram_s_38_2(ram_s_38_2), .n1193(n1193), .ram_s_38_1(ram_s_38_1), 
          .n1192(n1192), .n1191(n1191), .n1190(n1190), .ram_s_37_6(ram_s_37_6), 
          .n1189(n1189), .ram_s_37_5(ram_s_37_5), .n1188(n1188), .ram_s_37_4(ram_s_37_4), 
          .n1187(n1187), .ram_s_37_3(ram_s_37_3), .n1186(n1186), .ram_s_37_2(ram_s_37_2), 
          .n1185(n1185), .ram_s_37_1(ram_s_37_1), .n1184(n1184), .n1183(n1183), 
          .n1182(n1182), .ram_s_36_6(ram_s_36_6), .n1181(n1181), .ram_s_36_5(ram_s_36_5), 
          .n1180(n1180), .ram_s_36_4(ram_s_36_4), .n1179(n1179), .ram_s_36_3(ram_s_36_3), 
          .n1178(n1178), .ram_s_36_2(ram_s_36_2), .n1177(n1177), .ram_s_36_1(ram_s_36_1), 
          .n1176(n1176), .n1175(n1175), .n1174(n1174), .ram_s_35_6(ram_s_35_6), 
          .n1173(n1173), .ram_s_35_5(ram_s_35_5), .n1172(n1172), .ram_s_35_4(ram_s_35_4), 
          .n1171(n1171), .ram_s_35_3(ram_s_35_3), .n1170(n1170), .n1169(n1169), 
          .n1168(n1168), .ram_s_35_0(ram_s_35_0), .n1167(n1167), .n1166(n1166), 
          .ram_s_34_6(ram_s_34_6), .n1165(n1165), .ram_s_34_5(ram_s_34_5), 
          .n1164(n1164), .ram_s_34_4(ram_s_34_4), .n1163(n1163), .ram_s_34_3(ram_s_34_3), 
          .n1162(n1162), .n1161(n1161), .n1160(n1160), .ram_s_34_0(ram_s_34_0), 
          .n1159(n1159), .n1158(n1158), .ram_s_33_6(ram_s_33_6), .n1157(n1157), 
          .ram_s_33_5(ram_s_33_5), .n1156(n1156), .ram_s_33_4(ram_s_33_4), 
          .n1155(n1155), .ram_s_33_3(ram_s_33_3), .n1154(n1154), .n1153(n1153), 
          .n1152(n1152), .ram_s_33_0(ram_s_33_0), .n1151(n1151), .n1150(n1150), 
          .ram_s_32_6(ram_s_32_6), .n1149(n1149), .ram_s_32_5(ram_s_32_5), 
          .n1148(n1148), .ram_s_32_4(ram_s_32_4), .n1147(n1147), .ram_s_32_3(ram_s_32_3), 
          .n1146(n1146), .n1145(n1145), .n1144(n1144), .ram_s_32_0(ram_s_32_0), 
          .n1051(n1051), .n1047(n1047), .n1046(n1046), .n1045(n1045), 
          .ram_s_0_2(ram_s_0_2), .n1044(n1044), .ram_s_12_3(ram_s_12_3), 
          .n1043(n1043), .n1042(n1042), .ram_s_11_1(ram_s_11_1), .n1041(n1041), 
          .n1040(n1040), .ram_s_12_1(ram_s_12_1), .n1038(n1038), .ram_s_11_4(ram_s_11_4), 
          .n182(n182), .n1037(n1037), .ram_s_12_4(ram_s_12_4), .n54(n54), 
          .n1036(n1036), .ram_s_11_7(ram_s_11_7), .n183(n183), .n1035(n1035), 
          .n55(n55), .n1034(n1034), .ram_s_12_7(ram_s_12_7), .n184(n184), 
          .n1033(n1033), .ram_s_12_2(ram_s_12_2), .n56(n56), .n1032(n1032), 
          .ram_s_11_5(ram_s_11_5), .n185(n185), .n1031(n1031), .n57(n57), 
          .n1030(n1030), .ram_s_12_0(ram_s_12_0), .n186(n186), .n1029(n1029), 
          .ram_s_11_3(ram_s_11_3), .n58(n58), .n187(n187), .n59(n59), 
          .n188(n188), .n60(n60), .n189(n189), .n61(n61), .n190(n190), 
          .n62(n62), .n191(n191), .n63(n63), .n192(n192), .n1017(n1017), 
          .ram_s_0_3(ram_s_0_3), .n64(n64), .n1016(n1016), .ram_s_0_4(ram_s_0_4), 
          .n193(n193), .n1015(n1015), .ram_s_0_5(ram_s_0_5), .n65(n65), 
          .n1014(n1014), .ram_s_0_6(ram_s_0_6), .n194(n194), .n1013(n1013), 
          .n66(n66), .n1012(n1012), .n195(n195), .n1011(n1011), .n67(n67), 
          .n1010(n1010), .ram_s_1_2(ram_s_1_2), .n1009(n1009), .ram_s_1_3(ram_s_1_3), 
          .n1008(n1008), .ram_s_1_4(ram_s_1_4), .n1007(n1007), .ram_s_1_5(ram_s_1_5), 
          .n1006(n1006), .ram_s_4_4(ram_s_4_4), .n1005(n1005), .n1004(n1004), 
          .n1003(n1003), .ram_s_5_0(ram_s_5_0), .n1002(n1002), .ram_s_4_6(ram_s_4_6), 
          .n1001(n1001), .ram_s_5_1(ram_s_5_1), .n998(n998), .ram_s_8_5(ram_s_8_5), 
          .n997(n997), .n996(n996), .n995(n995), .ram_s_7_4(ram_s_7_4), 
          .n994(n994), .ram_s_7_1(ram_s_7_1), .n993(n993), .ram_s_6_6(ram_s_6_6), 
          .n992(n992), .ram_s_6_3(ram_s_6_3), .n989(n989), .n988(n988), 
          .ram_s_8_3(ram_s_8_3), .n987(n987), .ram_s_8_0(ram_s_8_0), .n986(n986), 
          .n199(n199), .n985(n985), .ram_s_7_2(ram_s_7_2), .n71(n71), 
          .n984(n984), .n200(n200), .n983(n983), .ram_s_6_4(ram_s_6_4), 
          .n72(n72), .n980(n980), .ram_s_8_7(ram_s_8_7), .n979(n979), 
          .ram_s_8_4(ram_s_8_4), .n978(n978), .ram_s_8_1(ram_s_8_1), .n977(n977), 
          .ram_s_7_6(ram_s_7_6), .n976(n976), .ram_s_7_3(ram_s_7_3), .n975(n975), 
          .ram_s_7_0(ram_s_7_0), .n974(n974), .n973(n973), .ram_s_1_6(ram_s_1_6), 
          .n972(n972), .n971(n971), .n970(n970), .n969(n969), .ram_s_2_2(ram_s_2_2), 
          .n968(n968), .ram_s_2_3(ram_s_2_3), .n967(n967), .ram_s_2_4(ram_s_2_4), 
          .n966(n966), .ram_s_2_5(ram_s_2_5), .n965(n965), .ram_s_2_6(ram_s_2_6), 
          .n964(n964), .n963(n963), .n962(n962), .n961(n961), .ram_s_3_2(ram_s_3_2), 
          .n960(n960), .ram_s_3_3(ram_s_3_3), .n959(n959), .ram_s_3_4(ram_s_3_4), 
          .n958(n958), .ram_s_3_5(ram_s_3_5), .n957(n957), .ram_s_14_7(ram_s_14_7), 
          .n952(n952), .ram_s_3_6(ram_s_3_6), .n950(n950), .n946(n946), 
          .ram_s_4_0(ram_s_4_0), .n944(n944), .ram_s_4_1(ram_s_4_1), .n941(n941), 
          .ram_s_4_2(ram_s_4_2), .n940(n940), .ram_s_5_2(ram_s_5_2), .n939(n939), 
          .ram_s_5_3(ram_s_5_3), .n935(n935), .n934(n934), .ram_s_6_0(ram_s_6_0), 
          .n933(n933), .ram_s_6_1(ram_s_6_1), .n932(n932), .ram_s_6_2(ram_s_6_2), 
          .n931(n931), .ram_s_5_6(ram_s_5_6), .n930(n930), .n927(n927), 
          .ram_s_4_3(ram_s_4_3), .n926(n926), .n925(n925), .ram_s_13_3(ram_s_13_3), 
          .n924(n924), .ram_s_13_4(ram_s_13_4), .n923(n923), .n210(n210), 
          .n82(n82), .n212(n212), .n84(n84), .n213(n213), .n85(n85), 
          .n214(n214), .n86(n86), .n217(n217), .n89(n89), .n218(n218), 
          .n90(n90), .n219(n219), .n91(n91), .n220(n220), .n92(n92), 
          .n221(n221), .n93(n93), .n222(n222), .n94(n94), .n223(n223), 
          .n95(n95), .n224(n224), .n96(n96), .n225(n225), .n97(n97), 
          .n918(n918), .ram_s_13_7(ram_s_13_7), .n917(n917), .ram_s_14_0(ram_s_14_0), 
          .n916(n916), .ram_s_14_1(ram_s_14_1), .n244(n244), .n116(n116), 
          .n115(n115), .n243(n243), .n245(n245), .n117(n117), .n246(n246), 
          .n118(n118), .n48(n48), .n176(n176), .n249(n249), .n121(n121), 
          .n250(n250), .n122(n122), .n251(n251), .n123(n123), .n252(n252), 
          .n124(n124), .n253(n253), .n125(n125), .n254(n254), .n126(n126), 
          .n255(n255), .n127(n127), .n256(n256), .n128(n128), .n257(n257), 
          .n129(n129), .ram_s_14_2(ram_s_14_2), .ram_s_13_2(ram_s_13_2), 
          .ram_s_11_0(ram_s_11_0), .n911(n911), .n909(n909), .n908(n908), 
          .ram_s_14_3(ram_s_14_3), .n907(n907), .ram_s_13_1(ram_s_13_1), 
          .n906(n906), .n904(n904), .ram_s_13_0(ram_s_13_0), .n901(n901), 
          .ram_s_5_4(ram_s_5_4), .n899(n899), .LED1_c_0(LED1_c_0), .n765(n765), 
          .n938(n938), .\pc_value[0] (pc_value[0]));   // src/top.vhd(96[23:28])
    SB_LUT4 i2312_3_lut (.I0(ram_s_209_0), .I1(register_vector[8]), .I2(n48), 
            .I3(GND_net), .O(n2560));   // src/ram.vhd(56[12:17])
    defparam i2312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2313_3_lut (.I0(ram_s_209_1), .I1(register_vector[9]), .I2(n48), 
            .I3(GND_net), .O(n2561));   // src/ram.vhd(56[12:17])
    defparam i2313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2314_3_lut (.I0(ram_s_209_2), .I1(register_vector[10]), .I2(n48), 
            .I3(GND_net), .O(n2562));   // src/ram.vhd(56[12:17])
    defparam i2314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2315_3_lut (.I0(ram_s_209_3), .I1(register_vector[11]), .I2(n48), 
            .I3(GND_net), .O(n2563));   // src/ram.vhd(56[12:17])
    defparam i2315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2316_3_lut (.I0(ram_s_209_4), .I1(sx[4]), .I2(n48), .I3(GND_net), 
            .O(n2564));   // src/ram.vhd(56[12:17])
    defparam i2316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2317_3_lut (.I0(ram_s_209_5), .I1(sx[5]), .I2(n48), .I3(GND_net), 
            .O(n2565));   // src/ram.vhd(56[12:17])
    defparam i2317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2318_3_lut (.I0(ram_s_209_6), .I1(sx[6]), .I2(n48), .I3(GND_net), 
            .O(n2566));   // src/ram.vhd(56[12:17])
    defparam i2318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1288_3_lut (.I0(ram_s_81_0), .I1(register_vector[8]), .I2(n176), 
            .I3(GND_net), .O(n1536));   // src/ram.vhd(56[12:17])
    defparam i1288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1289_3_lut (.I0(ram_s_81_1), .I1(register_vector[9]), .I2(n176), 
            .I3(GND_net), .O(n1537));   // src/ram.vhd(56[12:17])
    defparam i1289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1290_3_lut (.I0(ram_s_81_2), .I1(register_vector[10]), .I2(n176), 
            .I3(GND_net), .O(n1538));   // src/ram.vhd(56[12:17])
    defparam i1290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2319_3_lut (.I0(ram_s_209_7), .I1(sx[7]), .I2(n48), .I3(GND_net), 
            .O(n2567));   // src/ram.vhd(56[12:17])
    defparam i2319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1291_3_lut (.I0(ram_s_81_3), .I1(register_vector[11]), .I2(n176), 
            .I3(GND_net), .O(n1539));   // src/ram.vhd(56[12:17])
    defparam i1291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1292_3_lut (.I0(ram_s_81_4), .I1(sx[4]), .I2(n176), .I3(GND_net), 
            .O(n1540));   // src/ram.vhd(56[12:17])
    defparam i1292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1293_3_lut (.I0(ram_s_81_5), .I1(sx[5]), .I2(n176), .I3(GND_net), 
            .O(n1541));   // src/ram.vhd(56[12:17])
    defparam i1293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1294_3_lut (.I0(ram_s_81_6), .I1(sx[6]), .I2(n176), .I3(GND_net), 
            .O(n1542));   // src/ram.vhd(56[12:17])
    defparam i1294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1295_3_lut (.I0(ram_s_81_7), .I1(sx[7]), .I2(n176), .I3(GND_net), 
            .O(n1543));   // src/ram.vhd(56[12:17])
    defparam i1295_3_lut.LUT_INIT = 16'hcaca;
    SB_GB_IO CLK_3P3_MHZ_pad (.PACKAGE_PIN(CLK_3P3_MHZ), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(CLK_3P3_MHZ_c));   // src/top.vhd(36[9:20])
    defparam CLK_3P3_MHZ_pad.PIN_TYPE = 6'b000001;
    defparam CLK_3P3_MHZ_pad.PULLUP = 1'b0;
    defparam CLK_3P3_MHZ_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_3P3_MHZ_pad.IO_STANDARD = "SB_LVCMOS";
    GND i1 (.Y(GND_net));
    SB_IO BTN1_pad (.PACKAGE_PIN(BTN1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(BTN1_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam BTN1_pad.PIN_TYPE = 6'b000001;
    defparam BTN1_pad.PULLUP = 1'b0;
    defparam BTN1_pad.NEG_TRIGGER = 1'b0;
    defparam BTN1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED1_pad (.PACKAGE_PIN(LED1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED1_c_0));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED1_pad.PIN_TYPE = 6'b011001;
    defparam LED1_pad.PULLUP = 1'b0;
    defparam LED1_pad.NEG_TRIGGER = 1'b0;
    defparam LED1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1664_3_lut (.I0(ram_s_128_0), .I1(register_vector[8]), .I2(n129), 
            .I3(GND_net), .O(n1912));   // src/ram.vhd(56[12:17])
    defparam i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1665_3_lut (.I0(ram_s_128_1), .I1(register_vector[9]), .I2(n129), 
            .I3(GND_net), .O(n1913));   // src/ram.vhd(56[12:17])
    defparam i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1666_3_lut (.I0(ram_s_128_2), .I1(register_vector[10]), .I2(n129), 
            .I3(GND_net), .O(n1914));   // src/ram.vhd(56[12:17])
    defparam i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1667_3_lut (.I0(ram_s_128_3), .I1(register_vector[11]), .I2(n129), 
            .I3(GND_net), .O(n1915));   // src/ram.vhd(56[12:17])
    defparam i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1668_3_lut (.I0(ram_s_128_4), .I1(sx[4]), .I2(n129), .I3(GND_net), 
            .O(n1916));   // src/ram.vhd(56[12:17])
    defparam i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1669_3_lut (.I0(ram_s_128_5), .I1(sx[5]), .I2(n129), .I3(GND_net), 
            .O(n1917));   // src/ram.vhd(56[12:17])
    defparam i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1670_3_lut (.I0(ram_s_128_6), .I1(sx[6]), .I2(n129), .I3(GND_net), 
            .O(n1918));   // src/ram.vhd(56[12:17])
    defparam i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1671_3_lut (.I0(ram_s_128_7), .I1(sx[7]), .I2(n129), .I3(GND_net), 
            .O(n1919));   // src/ram.vhd(56[12:17])
    defparam i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1672_3_lut (.I0(ram_s_129_0), .I1(register_vector[8]), .I2(n128), 
            .I3(GND_net), .O(n1920));   // src/ram.vhd(56[12:17])
    defparam i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1673_3_lut (.I0(ram_s_129_1), .I1(register_vector[9]), .I2(n128), 
            .I3(GND_net), .O(n1921));   // src/ram.vhd(56[12:17])
    defparam i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1674_3_lut (.I0(ram_s_129_2), .I1(register_vector[10]), .I2(n128), 
            .I3(GND_net), .O(n1922));   // src/ram.vhd(56[12:17])
    defparam i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1675_3_lut (.I0(ram_s_129_3), .I1(register_vector[11]), .I2(n128), 
            .I3(GND_net), .O(n1923));   // src/ram.vhd(56[12:17])
    defparam i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1676_3_lut (.I0(ram_s_129_4), .I1(sx[4]), .I2(n128), .I3(GND_net), 
            .O(n1924));   // src/ram.vhd(56[12:17])
    defparam i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1677_3_lut (.I0(ram_s_129_5), .I1(sx[5]), .I2(n128), .I3(GND_net), 
            .O(n1925));   // src/ram.vhd(56[12:17])
    defparam i1677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1678_3_lut (.I0(ram_s_129_6), .I1(sx[6]), .I2(n128), .I3(GND_net), 
            .O(n1926));   // src/ram.vhd(56[12:17])
    defparam i1678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1679_3_lut (.I0(ram_s_129_7), .I1(sx[7]), .I2(n128), .I3(GND_net), 
            .O(n1927));   // src/ram.vhd(56[12:17])
    defparam i1679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1680_3_lut (.I0(ram_s_130_0), .I1(register_vector[8]), .I2(n127), 
            .I3(GND_net), .O(n1928));   // src/ram.vhd(56[12:17])
    defparam i1680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1681_3_lut (.I0(ram_s_130_1), .I1(register_vector[9]), .I2(n127), 
            .I3(GND_net), .O(n1929));   // src/ram.vhd(56[12:17])
    defparam i1681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1682_3_lut (.I0(ram_s_130_2), .I1(register_vector[10]), .I2(n127), 
            .I3(GND_net), .O(n1930));   // src/ram.vhd(56[12:17])
    defparam i1682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1683_3_lut (.I0(ram_s_130_3), .I1(register_vector[11]), .I2(n127), 
            .I3(GND_net), .O(n1931));   // src/ram.vhd(56[12:17])
    defparam i1683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1684_3_lut (.I0(ram_s_130_4), .I1(sx[4]), .I2(n127), .I3(GND_net), 
            .O(n1932));   // src/ram.vhd(56[12:17])
    defparam i1684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1685_3_lut (.I0(ram_s_130_5), .I1(sx[5]), .I2(n127), .I3(GND_net), 
            .O(n1933));   // src/ram.vhd(56[12:17])
    defparam i1685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1686_3_lut (.I0(ram_s_130_6), .I1(sx[6]), .I2(n127), .I3(GND_net), 
            .O(n1934));   // src/ram.vhd(56[12:17])
    defparam i1686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1687_3_lut (.I0(ram_s_130_7), .I1(sx[7]), .I2(n127), .I3(GND_net), 
            .O(n1935));   // src/ram.vhd(56[12:17])
    defparam i1687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1688_3_lut (.I0(ram_s_131_0), .I1(register_vector[8]), .I2(n126), 
            .I3(GND_net), .O(n1936));   // src/ram.vhd(56[12:17])
    defparam i1688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1689_3_lut (.I0(ram_s_131_1), .I1(register_vector[9]), .I2(n126), 
            .I3(GND_net), .O(n1937));   // src/ram.vhd(56[12:17])
    defparam i1689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1690_3_lut (.I0(ram_s_131_2), .I1(register_vector[10]), .I2(n126), 
            .I3(GND_net), .O(n1938));   // src/ram.vhd(56[12:17])
    defparam i1690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1691_3_lut (.I0(ram_s_131_3), .I1(register_vector[11]), .I2(n126), 
            .I3(GND_net), .O(n1939));   // src/ram.vhd(56[12:17])
    defparam i1691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1692_3_lut (.I0(ram_s_131_4), .I1(sx[4]), .I2(n126), .I3(GND_net), 
            .O(n1940));   // src/ram.vhd(56[12:17])
    defparam i1692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1693_3_lut (.I0(ram_s_131_5), .I1(sx[5]), .I2(n126), .I3(GND_net), 
            .O(n1941));   // src/ram.vhd(56[12:17])
    defparam i1693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1694_3_lut (.I0(ram_s_131_6), .I1(sx[6]), .I2(n126), .I3(GND_net), 
            .O(n1942));   // src/ram.vhd(56[12:17])
    defparam i1694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1695_3_lut (.I0(ram_s_131_7), .I1(sx[7]), .I2(n126), .I3(GND_net), 
            .O(n1943));   // src/ram.vhd(56[12:17])
    defparam i1695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1696_3_lut (.I0(ram_s_132_0), .I1(register_vector[8]), .I2(n125), 
            .I3(GND_net), .O(n1944));   // src/ram.vhd(56[12:17])
    defparam i1696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1697_3_lut (.I0(ram_s_132_1), .I1(register_vector[9]), .I2(n125), 
            .I3(GND_net), .O(n1945));   // src/ram.vhd(56[12:17])
    defparam i1697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1698_3_lut (.I0(ram_s_132_2), .I1(register_vector[10]), .I2(n125), 
            .I3(GND_net), .O(n1946));   // src/ram.vhd(56[12:17])
    defparam i1698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1699_3_lut (.I0(ram_s_132_3), .I1(register_vector[11]), .I2(n125), 
            .I3(GND_net), .O(n1947));   // src/ram.vhd(56[12:17])
    defparam i1699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1700_3_lut (.I0(ram_s_132_4), .I1(sx[4]), .I2(n125), .I3(GND_net), 
            .O(n1948));   // src/ram.vhd(56[12:17])
    defparam i1700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1701_3_lut (.I0(ram_s_132_5), .I1(sx[5]), .I2(n125), .I3(GND_net), 
            .O(n1949));   // src/ram.vhd(56[12:17])
    defparam i1701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1702_3_lut (.I0(ram_s_132_6), .I1(sx[6]), .I2(n125), .I3(GND_net), 
            .O(n1950));   // src/ram.vhd(56[12:17])
    defparam i1702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1703_3_lut (.I0(ram_s_132_7), .I1(sx[7]), .I2(n125), .I3(GND_net), 
            .O(n1951));   // src/ram.vhd(56[12:17])
    defparam i1703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1704_3_lut (.I0(ram_s_133_0), .I1(register_vector[8]), .I2(n124), 
            .I3(GND_net), .O(n1952));   // src/ram.vhd(56[12:17])
    defparam i1704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1705_3_lut (.I0(ram_s_133_1), .I1(register_vector[9]), .I2(n124), 
            .I3(GND_net), .O(n1953));   // src/ram.vhd(56[12:17])
    defparam i1705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1706_3_lut (.I0(ram_s_133_2), .I1(register_vector[10]), .I2(n124), 
            .I3(GND_net), .O(n1954));   // src/ram.vhd(56[12:17])
    defparam i1706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1707_3_lut (.I0(ram_s_133_3), .I1(register_vector[11]), .I2(n124), 
            .I3(GND_net), .O(n1955));   // src/ram.vhd(56[12:17])
    defparam i1707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1708_3_lut (.I0(ram_s_133_4), .I1(sx[4]), .I2(n124), .I3(GND_net), 
            .O(n1956));   // src/ram.vhd(56[12:17])
    defparam i1708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1709_3_lut (.I0(ram_s_133_5), .I1(sx[5]), .I2(n124), .I3(GND_net), 
            .O(n1957));   // src/ram.vhd(56[12:17])
    defparam i1709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1710_3_lut (.I0(ram_s_133_6), .I1(sx[6]), .I2(n124), .I3(GND_net), 
            .O(n1958));   // src/ram.vhd(56[12:17])
    defparam i1710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1711_3_lut (.I0(ram_s_133_7), .I1(sx[7]), .I2(n124), .I3(GND_net), 
            .O(n1959));   // src/ram.vhd(56[12:17])
    defparam i1711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1712_3_lut (.I0(ram_s_134_0), .I1(register_vector[8]), .I2(n123), 
            .I3(GND_net), .O(n1960));   // src/ram.vhd(56[12:17])
    defparam i1712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1713_3_lut (.I0(ram_s_134_1), .I1(register_vector[9]), .I2(n123), 
            .I3(GND_net), .O(n1961));   // src/ram.vhd(56[12:17])
    defparam i1713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1714_3_lut (.I0(ram_s_134_2), .I1(register_vector[10]), .I2(n123), 
            .I3(GND_net), .O(n1962));   // src/ram.vhd(56[12:17])
    defparam i1714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1715_3_lut (.I0(ram_s_134_3), .I1(register_vector[11]), .I2(n123), 
            .I3(GND_net), .O(n1963));   // src/ram.vhd(56[12:17])
    defparam i1715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1716_3_lut (.I0(ram_s_134_4), .I1(sx[4]), .I2(n123), .I3(GND_net), 
            .O(n1964));   // src/ram.vhd(56[12:17])
    defparam i1716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1717_3_lut (.I0(ram_s_134_5), .I1(sx[5]), .I2(n123), .I3(GND_net), 
            .O(n1965));   // src/ram.vhd(56[12:17])
    defparam i1717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1718_3_lut (.I0(ram_s_134_6), .I1(sx[6]), .I2(n123), .I3(GND_net), 
            .O(n1966));   // src/ram.vhd(56[12:17])
    defparam i1718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1719_3_lut (.I0(ram_s_134_7), .I1(sx[7]), .I2(n123), .I3(GND_net), 
            .O(n1967));   // src/ram.vhd(56[12:17])
    defparam i1719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1720_3_lut (.I0(ram_s_135_0), .I1(register_vector[8]), .I2(n122), 
            .I3(GND_net), .O(n1968));   // src/ram.vhd(56[12:17])
    defparam i1720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1721_3_lut (.I0(ram_s_135_1), .I1(register_vector[9]), .I2(n122), 
            .I3(GND_net), .O(n1969));   // src/ram.vhd(56[12:17])
    defparam i1721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1722_3_lut (.I0(ram_s_135_2), .I1(register_vector[10]), .I2(n122), 
            .I3(GND_net), .O(n1970));   // src/ram.vhd(56[12:17])
    defparam i1722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1723_3_lut (.I0(ram_s_135_3), .I1(register_vector[11]), .I2(n122), 
            .I3(GND_net), .O(n1971));   // src/ram.vhd(56[12:17])
    defparam i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1724_3_lut (.I0(ram_s_135_4), .I1(sx[4]), .I2(n122), .I3(GND_net), 
            .O(n1972));   // src/ram.vhd(56[12:17])
    defparam i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1725_3_lut (.I0(ram_s_135_5), .I1(sx[5]), .I2(n122), .I3(GND_net), 
            .O(n1973));   // src/ram.vhd(56[12:17])
    defparam i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1726_3_lut (.I0(ram_s_135_6), .I1(sx[6]), .I2(n122), .I3(GND_net), 
            .O(n1974));   // src/ram.vhd(56[12:17])
    defparam i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1727_3_lut (.I0(ram_s_135_7), .I1(sx[7]), .I2(n122), .I3(GND_net), 
            .O(n1975));   // src/ram.vhd(56[12:17])
    defparam i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1728_3_lut (.I0(ram_s_136_0), .I1(register_vector[8]), .I2(n121), 
            .I3(GND_net), .O(n1976));   // src/ram.vhd(56[12:17])
    defparam i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1729_3_lut (.I0(ram_s_136_1), .I1(register_vector[9]), .I2(n121), 
            .I3(GND_net), .O(n1977));   // src/ram.vhd(56[12:17])
    defparam i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1730_3_lut (.I0(ram_s_136_2), .I1(register_vector[10]), .I2(n121), 
            .I3(GND_net), .O(n1978));   // src/ram.vhd(56[12:17])
    defparam i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1731_3_lut (.I0(ram_s_136_3), .I1(register_vector[11]), .I2(n121), 
            .I3(GND_net), .O(n1979));   // src/ram.vhd(56[12:17])
    defparam i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1732_3_lut (.I0(ram_s_136_4), .I1(sx[4]), .I2(n121), .I3(GND_net), 
            .O(n1980));   // src/ram.vhd(56[12:17])
    defparam i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1733_3_lut (.I0(ram_s_136_5), .I1(sx[5]), .I2(n121), .I3(GND_net), 
            .O(n1981));   // src/ram.vhd(56[12:17])
    defparam i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1734_3_lut (.I0(ram_s_136_6), .I1(sx[6]), .I2(n121), .I3(GND_net), 
            .O(n1982));   // src/ram.vhd(56[12:17])
    defparam i1734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1735_3_lut (.I0(ram_s_136_7), .I1(sx[7]), .I2(n121), .I3(GND_net), 
            .O(n1983));   // src/ram.vhd(56[12:17])
    defparam i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1752_3_lut (.I0(ram_s_139_0), .I1(register_vector[8]), .I2(n118), 
            .I3(GND_net), .O(n2000));   // src/ram.vhd(56[12:17])
    defparam i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1753_3_lut (.I0(ram_s_139_1), .I1(register_vector[9]), .I2(n118), 
            .I3(GND_net), .O(n2001));   // src/ram.vhd(56[12:17])
    defparam i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1754_3_lut (.I0(ram_s_139_2), .I1(register_vector[10]), .I2(n118), 
            .I3(GND_net), .O(n2002));   // src/ram.vhd(56[12:17])
    defparam i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1755_3_lut (.I0(ram_s_139_3), .I1(register_vector[11]), .I2(n118), 
            .I3(GND_net), .O(n2003));   // src/ram.vhd(56[12:17])
    defparam i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1756_3_lut (.I0(ram_s_139_4), .I1(sx[4]), .I2(n118), .I3(GND_net), 
            .O(n2004));   // src/ram.vhd(56[12:17])
    defparam i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1757_3_lut (.I0(ram_s_139_5), .I1(sx[5]), .I2(n118), .I3(GND_net), 
            .O(n2005));   // src/ram.vhd(56[12:17])
    defparam i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1758_3_lut (.I0(ram_s_139_6), .I1(sx[6]), .I2(n118), .I3(GND_net), 
            .O(n2006));   // src/ram.vhd(56[12:17])
    defparam i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1759_3_lut (.I0(ram_s_139_7), .I1(sx[7]), .I2(n118), .I3(GND_net), 
            .O(n2007));   // src/ram.vhd(56[12:17])
    defparam i1759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1760_3_lut (.I0(ram_s_140_0), .I1(register_vector[8]), .I2(n117), 
            .I3(GND_net), .O(n2008));   // src/ram.vhd(56[12:17])
    defparam i1760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1761_3_lut (.I0(ram_s_140_1), .I1(register_vector[9]), .I2(n117), 
            .I3(GND_net), .O(n2009));   // src/ram.vhd(56[12:17])
    defparam i1761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1762_3_lut (.I0(ram_s_140_2), .I1(register_vector[10]), .I2(n117), 
            .I3(GND_net), .O(n2010));   // src/ram.vhd(56[12:17])
    defparam i1762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1763_3_lut (.I0(ram_s_140_3), .I1(register_vector[11]), .I2(n117), 
            .I3(GND_net), .O(n2011));   // src/ram.vhd(56[12:17])
    defparam i1763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1764_3_lut (.I0(ram_s_140_4), .I1(sx[4]), .I2(n117), .I3(GND_net), 
            .O(n2012));   // src/ram.vhd(56[12:17])
    defparam i1764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1765_3_lut (.I0(ram_s_140_5), .I1(sx[5]), .I2(n117), .I3(GND_net), 
            .O(n2013));   // src/ram.vhd(56[12:17])
    defparam i1765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1766_3_lut (.I0(ram_s_140_6), .I1(sx[6]), .I2(n117), .I3(GND_net), 
            .O(n2014));   // src/ram.vhd(56[12:17])
    defparam i1766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1767_3_lut (.I0(ram_s_140_7), .I1(sx[7]), .I2(n117), .I3(GND_net), 
            .O(n2015));   // src/ram.vhd(56[12:17])
    defparam i1767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i645_3_lut (.I0(ram_s_14_4), .I1(sx[4]), .I2(n243), .I3(GND_net), 
            .O(n893));   // src/ram.vhd(56[12:17])
    defparam i645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1768_3_lut (.I0(ram_s_141_0), .I1(register_vector[8]), .I2(n116), 
            .I3(GND_net), .O(n2016));   // src/ram.vhd(56[12:17])
    defparam i1768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1769_3_lut (.I0(ram_s_141_1), .I1(register_vector[9]), .I2(n116), 
            .I3(GND_net), .O(n2017));   // src/ram.vhd(56[12:17])
    defparam i1769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1770_3_lut (.I0(ram_s_141_2), .I1(register_vector[10]), .I2(n116), 
            .I3(GND_net), .O(n2018));   // src/ram.vhd(56[12:17])
    defparam i1770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1771_3_lut (.I0(ram_s_141_3), .I1(register_vector[11]), .I2(n116), 
            .I3(GND_net), .O(n2019));   // src/ram.vhd(56[12:17])
    defparam i1771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1772_3_lut (.I0(ram_s_141_4), .I1(sx[4]), .I2(n116), .I3(GND_net), 
            .O(n2020));   // src/ram.vhd(56[12:17])
    defparam i1772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1773_3_lut (.I0(ram_s_141_5), .I1(sx[5]), .I2(n116), .I3(GND_net), 
            .O(n2021));   // src/ram.vhd(56[12:17])
    defparam i1773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1774_3_lut (.I0(ram_s_141_6), .I1(sx[6]), .I2(n116), .I3(GND_net), 
            .O(n2022));   // src/ram.vhd(56[12:17])
    defparam i1774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1775_3_lut (.I0(ram_s_141_7), .I1(sx[7]), .I2(n116), .I3(GND_net), 
            .O(n2023));   // src/ram.vhd(56[12:17])
    defparam i1775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1776_3_lut (.I0(ram_s_142_0), .I1(register_vector[8]), .I2(n115), 
            .I3(GND_net), .O(n2024));   // src/ram.vhd(56[12:17])
    defparam i1776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1777_3_lut (.I0(ram_s_142_1), .I1(register_vector[9]), .I2(n115), 
            .I3(GND_net), .O(n2025));   // src/ram.vhd(56[12:17])
    defparam i1777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1778_3_lut (.I0(ram_s_142_2), .I1(register_vector[10]), .I2(n115), 
            .I3(GND_net), .O(n2026));   // src/ram.vhd(56[12:17])
    defparam i1778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1779_3_lut (.I0(ram_s_142_3), .I1(register_vector[11]), .I2(n115), 
            .I3(GND_net), .O(n2027));   // src/ram.vhd(56[12:17])
    defparam i1779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1780_3_lut (.I0(ram_s_142_4), .I1(sx[4]), .I2(n115), .I3(GND_net), 
            .O(n2028));   // src/ram.vhd(56[12:17])
    defparam i1780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1781_3_lut (.I0(ram_s_142_5), .I1(sx[5]), .I2(n115), .I3(GND_net), 
            .O(n2029));   // src/ram.vhd(56[12:17])
    defparam i1781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1782_3_lut (.I0(ram_s_142_6), .I1(sx[6]), .I2(n115), .I3(GND_net), 
            .O(n2030));   // src/ram.vhd(56[12:17])
    defparam i1782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1783_3_lut (.I0(ram_s_142_7), .I1(sx[7]), .I2(n115), .I3(GND_net), 
            .O(n2031));   // src/ram.vhd(56[12:17])
    defparam i1783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(internal_reset), .I1(special_bit), .I2(bram_enable), 
            .I3(t_state[1]), .O(n8580));   // src/state_machine.vhd(70[9] 79[16])
    defparam i1_4_lut.LUT_INIT = 16'h1505;
    SB_LUT4 i1_2_lut (.I0(t_state[1]), .I1(internal_reset), .I2(GND_net), 
            .I3(GND_net), .O(n765));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1920_3_lut (.I0(ram_s_160_0), .I1(register_vector[8]), .I2(n97), 
            .I3(GND_net), .O(n2168));   // src/ram.vhd(56[12:17])
    defparam i1920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1921_3_lut (.I0(ram_s_160_1), .I1(register_vector[9]), .I2(n97), 
            .I3(GND_net), .O(n2169));   // src/ram.vhd(56[12:17])
    defparam i1921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1922_3_lut (.I0(ram_s_160_2), .I1(register_vector[10]), .I2(n97), 
            .I3(GND_net), .O(n2170));   // src/ram.vhd(56[12:17])
    defparam i1922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1923_3_lut (.I0(ram_s_160_3), .I1(register_vector[11]), .I2(n97), 
            .I3(GND_net), .O(n2171));   // src/ram.vhd(56[12:17])
    defparam i1923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1924_3_lut (.I0(ram_s_160_4), .I1(sx[4]), .I2(n97), .I3(GND_net), 
            .O(n2172));   // src/ram.vhd(56[12:17])
    defparam i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1925_3_lut (.I0(ram_s_160_5), .I1(sx[5]), .I2(n97), .I3(GND_net), 
            .O(n2173));   // src/ram.vhd(56[12:17])
    defparam i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1926_3_lut (.I0(ram_s_160_6), .I1(sx[6]), .I2(n97), .I3(GND_net), 
            .O(n2174));   // src/ram.vhd(56[12:17])
    defparam i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1927_3_lut (.I0(ram_s_160_7), .I1(sx[7]), .I2(n97), .I3(GND_net), 
            .O(n2175));   // src/ram.vhd(56[12:17])
    defparam i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1928_3_lut (.I0(ram_s_161_0), .I1(register_vector[8]), .I2(n96), 
            .I3(GND_net), .O(n2176));   // src/ram.vhd(56[12:17])
    defparam i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1929_3_lut (.I0(ram_s_161_1), .I1(register_vector[9]), .I2(n96), 
            .I3(GND_net), .O(n2177));   // src/ram.vhd(56[12:17])
    defparam i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1930_3_lut (.I0(ram_s_161_2), .I1(register_vector[10]), .I2(n96), 
            .I3(GND_net), .O(n2178));   // src/ram.vhd(56[12:17])
    defparam i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1931_3_lut (.I0(ram_s_161_3), .I1(register_vector[11]), .I2(n96), 
            .I3(GND_net), .O(n2179));   // src/ram.vhd(56[12:17])
    defparam i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1932_3_lut (.I0(ram_s_161_4), .I1(sx[4]), .I2(n96), .I3(GND_net), 
            .O(n2180));   // src/ram.vhd(56[12:17])
    defparam i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1933_3_lut (.I0(ram_s_161_5), .I1(sx[5]), .I2(n96), .I3(GND_net), 
            .O(n2181));   // src/ram.vhd(56[12:17])
    defparam i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1934_3_lut (.I0(ram_s_161_6), .I1(sx[6]), .I2(n96), .I3(GND_net), 
            .O(n2182));   // src/ram.vhd(56[12:17])
    defparam i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1935_3_lut (.I0(ram_s_161_7), .I1(sx[7]), .I2(n96), .I3(GND_net), 
            .O(n2183));   // src/ram.vhd(56[12:17])
    defparam i1935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1936_3_lut (.I0(ram_s_162_0), .I1(register_vector[8]), .I2(n95), 
            .I3(GND_net), .O(n2184));   // src/ram.vhd(56[12:17])
    defparam i1936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1937_3_lut (.I0(ram_s_162_1), .I1(register_vector[9]), .I2(n95), 
            .I3(GND_net), .O(n2185));   // src/ram.vhd(56[12:17])
    defparam i1937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1938_3_lut (.I0(ram_s_162_2), .I1(register_vector[10]), .I2(n95), 
            .I3(GND_net), .O(n2186));   // src/ram.vhd(56[12:17])
    defparam i1938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1939_3_lut (.I0(ram_s_162_3), .I1(register_vector[11]), .I2(n95), 
            .I3(GND_net), .O(n2187));   // src/ram.vhd(56[12:17])
    defparam i1939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1940_3_lut (.I0(ram_s_162_4), .I1(sx[4]), .I2(n95), .I3(GND_net), 
            .O(n2188));   // src/ram.vhd(56[12:17])
    defparam i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1941_3_lut (.I0(ram_s_162_5), .I1(sx[5]), .I2(n95), .I3(GND_net), 
            .O(n2189));   // src/ram.vhd(56[12:17])
    defparam i1941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1942_3_lut (.I0(ram_s_162_6), .I1(sx[6]), .I2(n95), .I3(GND_net), 
            .O(n2190));   // src/ram.vhd(56[12:17])
    defparam i1942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1943_3_lut (.I0(ram_s_162_7), .I1(sx[7]), .I2(n95), .I3(GND_net), 
            .O(n2191));   // src/ram.vhd(56[12:17])
    defparam i1943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1944_3_lut (.I0(ram_s_163_0), .I1(register_vector[8]), .I2(n94), 
            .I3(GND_net), .O(n2192));   // src/ram.vhd(56[12:17])
    defparam i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1945_3_lut (.I0(ram_s_163_1), .I1(register_vector[9]), .I2(n94), 
            .I3(GND_net), .O(n2193));   // src/ram.vhd(56[12:17])
    defparam i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1946_3_lut (.I0(ram_s_163_2), .I1(register_vector[10]), .I2(n94), 
            .I3(GND_net), .O(n2194));   // src/ram.vhd(56[12:17])
    defparam i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1947_3_lut (.I0(ram_s_163_3), .I1(register_vector[11]), .I2(n94), 
            .I3(GND_net), .O(n2195));   // src/ram.vhd(56[12:17])
    defparam i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1948_3_lut (.I0(ram_s_163_4), .I1(sx[4]), .I2(n94), .I3(GND_net), 
            .O(n2196));   // src/ram.vhd(56[12:17])
    defparam i1948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1949_3_lut (.I0(ram_s_163_5), .I1(sx[5]), .I2(n94), .I3(GND_net), 
            .O(n2197));   // src/ram.vhd(56[12:17])
    defparam i1949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1950_3_lut (.I0(ram_s_163_6), .I1(sx[6]), .I2(n94), .I3(GND_net), 
            .O(n2198));   // src/ram.vhd(56[12:17])
    defparam i1950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1951_3_lut (.I0(ram_s_163_7), .I1(sx[7]), .I2(n94), .I3(GND_net), 
            .O(n2199));   // src/ram.vhd(56[12:17])
    defparam i1951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1952_3_lut (.I0(ram_s_164_0), .I1(register_vector[8]), .I2(n93), 
            .I3(GND_net), .O(n2200));   // src/ram.vhd(56[12:17])
    defparam i1952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1953_3_lut (.I0(ram_s_164_1), .I1(register_vector[9]), .I2(n93), 
            .I3(GND_net), .O(n2201));   // src/ram.vhd(56[12:17])
    defparam i1953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1954_3_lut (.I0(ram_s_164_2), .I1(register_vector[10]), .I2(n93), 
            .I3(GND_net), .O(n2202));   // src/ram.vhd(56[12:17])
    defparam i1954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1955_3_lut (.I0(ram_s_164_3), .I1(register_vector[11]), .I2(n93), 
            .I3(GND_net), .O(n2203));   // src/ram.vhd(56[12:17])
    defparam i1955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1956_3_lut (.I0(ram_s_164_4), .I1(sx[4]), .I2(n93), .I3(GND_net), 
            .O(n2204));   // src/ram.vhd(56[12:17])
    defparam i1956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1957_3_lut (.I0(ram_s_164_5), .I1(sx[5]), .I2(n93), .I3(GND_net), 
            .O(n2205));   // src/ram.vhd(56[12:17])
    defparam i1957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1958_3_lut (.I0(ram_s_164_6), .I1(sx[6]), .I2(n93), .I3(GND_net), 
            .O(n2206));   // src/ram.vhd(56[12:17])
    defparam i1958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1959_3_lut (.I0(ram_s_164_7), .I1(sx[7]), .I2(n93), .I3(GND_net), 
            .O(n2207));   // src/ram.vhd(56[12:17])
    defparam i1959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1960_3_lut (.I0(ram_s_165_0), .I1(register_vector[8]), .I2(n92), 
            .I3(GND_net), .O(n2208));   // src/ram.vhd(56[12:17])
    defparam i1960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1961_3_lut (.I0(ram_s_165_1), .I1(register_vector[9]), .I2(n92), 
            .I3(GND_net), .O(n2209));   // src/ram.vhd(56[12:17])
    defparam i1961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1962_3_lut (.I0(ram_s_165_2), .I1(register_vector[10]), .I2(n92), 
            .I3(GND_net), .O(n2210));   // src/ram.vhd(56[12:17])
    defparam i1962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1963_3_lut (.I0(ram_s_165_3), .I1(register_vector[11]), .I2(n92), 
            .I3(GND_net), .O(n2211));   // src/ram.vhd(56[12:17])
    defparam i1963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1964_3_lut (.I0(ram_s_165_4), .I1(sx[4]), .I2(n92), .I3(GND_net), 
            .O(n2212));   // src/ram.vhd(56[12:17])
    defparam i1964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1965_3_lut (.I0(ram_s_165_5), .I1(sx[5]), .I2(n92), .I3(GND_net), 
            .O(n2213));   // src/ram.vhd(56[12:17])
    defparam i1965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1966_3_lut (.I0(ram_s_165_6), .I1(sx[6]), .I2(n92), .I3(GND_net), 
            .O(n2214));   // src/ram.vhd(56[12:17])
    defparam i1966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1967_3_lut (.I0(ram_s_165_7), .I1(sx[7]), .I2(n92), .I3(GND_net), 
            .O(n2215));   // src/ram.vhd(56[12:17])
    defparam i1967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1968_3_lut (.I0(ram_s_166_0), .I1(register_vector[8]), .I2(n91), 
            .I3(GND_net), .O(n2216));   // src/ram.vhd(56[12:17])
    defparam i1968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1969_3_lut (.I0(ram_s_166_1), .I1(register_vector[9]), .I2(n91), 
            .I3(GND_net), .O(n2217));   // src/ram.vhd(56[12:17])
    defparam i1969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1970_3_lut (.I0(ram_s_166_2), .I1(register_vector[10]), .I2(n91), 
            .I3(GND_net), .O(n2218));   // src/ram.vhd(56[12:17])
    defparam i1970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1971_3_lut (.I0(ram_s_166_3), .I1(register_vector[11]), .I2(n91), 
            .I3(GND_net), .O(n2219));   // src/ram.vhd(56[12:17])
    defparam i1971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1972_3_lut (.I0(ram_s_166_4), .I1(sx[4]), .I2(n91), .I3(GND_net), 
            .O(n2220));   // src/ram.vhd(56[12:17])
    defparam i1972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1973_3_lut (.I0(ram_s_166_5), .I1(sx[5]), .I2(n91), .I3(GND_net), 
            .O(n2221));   // src/ram.vhd(56[12:17])
    defparam i1973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1974_3_lut (.I0(ram_s_166_6), .I1(sx[6]), .I2(n91), .I3(GND_net), 
            .O(n2222));   // src/ram.vhd(56[12:17])
    defparam i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1975_3_lut (.I0(ram_s_166_7), .I1(sx[7]), .I2(n91), .I3(GND_net), 
            .O(n2223));   // src/ram.vhd(56[12:17])
    defparam i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1976_3_lut (.I0(ram_s_167_0), .I1(register_vector[8]), .I2(n90), 
            .I3(GND_net), .O(n2224));   // src/ram.vhd(56[12:17])
    defparam i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1977_3_lut (.I0(ram_s_167_1), .I1(register_vector[9]), .I2(n90), 
            .I3(GND_net), .O(n2225));   // src/ram.vhd(56[12:17])
    defparam i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1978_3_lut (.I0(ram_s_167_2), .I1(register_vector[10]), .I2(n90), 
            .I3(GND_net), .O(n2226));   // src/ram.vhd(56[12:17])
    defparam i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1979_3_lut (.I0(ram_s_167_3), .I1(register_vector[11]), .I2(n90), 
            .I3(GND_net), .O(n2227));   // src/ram.vhd(56[12:17])
    defparam i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1980_3_lut (.I0(ram_s_167_4), .I1(sx[4]), .I2(n90), .I3(GND_net), 
            .O(n2228));   // src/ram.vhd(56[12:17])
    defparam i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1981_3_lut (.I0(ram_s_167_5), .I1(sx[5]), .I2(n90), .I3(GND_net), 
            .O(n2229));   // src/ram.vhd(56[12:17])
    defparam i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1982_3_lut (.I0(ram_s_167_6), .I1(sx[6]), .I2(n90), .I3(GND_net), 
            .O(n2230));   // src/ram.vhd(56[12:17])
    defparam i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1983_3_lut (.I0(ram_s_167_7), .I1(sx[7]), .I2(n90), .I3(GND_net), 
            .O(n2231));   // src/ram.vhd(56[12:17])
    defparam i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1984_3_lut (.I0(ram_s_168_0), .I1(register_vector[8]), .I2(n89), 
            .I3(GND_net), .O(n2232));   // src/ram.vhd(56[12:17])
    defparam i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1985_3_lut (.I0(ram_s_168_1), .I1(register_vector[9]), .I2(n89), 
            .I3(GND_net), .O(n2233));   // src/ram.vhd(56[12:17])
    defparam i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1986_3_lut (.I0(ram_s_168_2), .I1(register_vector[10]), .I2(n89), 
            .I3(GND_net), .O(n2234));   // src/ram.vhd(56[12:17])
    defparam i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1987_3_lut (.I0(ram_s_168_3), .I1(register_vector[11]), .I2(n89), 
            .I3(GND_net), .O(n2235));   // src/ram.vhd(56[12:17])
    defparam i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1988_3_lut (.I0(ram_s_168_4), .I1(sx[4]), .I2(n89), .I3(GND_net), 
            .O(n2236));   // src/ram.vhd(56[12:17])
    defparam i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1989_3_lut (.I0(ram_s_168_5), .I1(sx[5]), .I2(n89), .I3(GND_net), 
            .O(n2237));   // src/ram.vhd(56[12:17])
    defparam i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1990_3_lut (.I0(ram_s_168_6), .I1(sx[6]), .I2(n89), .I3(GND_net), 
            .O(n2238));   // src/ram.vhd(56[12:17])
    defparam i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1991_3_lut (.I0(ram_s_168_7), .I1(sx[7]), .I2(n89), .I3(GND_net), 
            .O(n2239));   // src/ram.vhd(56[12:17])
    defparam i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2008_3_lut (.I0(ram_s_171_0), .I1(register_vector[8]), .I2(n86), 
            .I3(GND_net), .O(n2256));   // src/ram.vhd(56[12:17])
    defparam i2008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2009_3_lut (.I0(ram_s_171_1), .I1(register_vector[9]), .I2(n86), 
            .I3(GND_net), .O(n2257));   // src/ram.vhd(56[12:17])
    defparam i2009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2010_3_lut (.I0(ram_s_171_2), .I1(register_vector[10]), .I2(n86), 
            .I3(GND_net), .O(n2258));   // src/ram.vhd(56[12:17])
    defparam i2010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2011_3_lut (.I0(ram_s_171_3), .I1(register_vector[11]), .I2(n86), 
            .I3(GND_net), .O(n2259));   // src/ram.vhd(56[12:17])
    defparam i2011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2012_3_lut (.I0(ram_s_171_4), .I1(sx[4]), .I2(n86), .I3(GND_net), 
            .O(n2260));   // src/ram.vhd(56[12:17])
    defparam i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2013_3_lut (.I0(ram_s_171_5), .I1(sx[5]), .I2(n86), .I3(GND_net), 
            .O(n2261));   // src/ram.vhd(56[12:17])
    defparam i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2014_3_lut (.I0(ram_s_171_6), .I1(sx[6]), .I2(n86), .I3(GND_net), 
            .O(n2262));   // src/ram.vhd(56[12:17])
    defparam i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2015_3_lut (.I0(ram_s_171_7), .I1(sx[7]), .I2(n86), .I3(GND_net), 
            .O(n2263));   // src/ram.vhd(56[12:17])
    defparam i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2016_3_lut (.I0(ram_s_172_0), .I1(register_vector[8]), .I2(n85), 
            .I3(GND_net), .O(n2264));   // src/ram.vhd(56[12:17])
    defparam i2016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2017_3_lut (.I0(ram_s_172_1), .I1(register_vector[9]), .I2(n85), 
            .I3(GND_net), .O(n2265));   // src/ram.vhd(56[12:17])
    defparam i2017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2018_3_lut (.I0(ram_s_172_2), .I1(register_vector[10]), .I2(n85), 
            .I3(GND_net), .O(n2266));   // src/ram.vhd(56[12:17])
    defparam i2018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2019_3_lut (.I0(ram_s_172_3), .I1(register_vector[11]), .I2(n85), 
            .I3(GND_net), .O(n2267));   // src/ram.vhd(56[12:17])
    defparam i2019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2020_3_lut (.I0(ram_s_172_4), .I1(sx[4]), .I2(n85), .I3(GND_net), 
            .O(n2268));   // src/ram.vhd(56[12:17])
    defparam i2020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2021_3_lut (.I0(ram_s_172_5), .I1(sx[5]), .I2(n85), .I3(GND_net), 
            .O(n2269));   // src/ram.vhd(56[12:17])
    defparam i2021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2022_3_lut (.I0(ram_s_172_6), .I1(sx[6]), .I2(n85), .I3(GND_net), 
            .O(n2270));   // src/ram.vhd(56[12:17])
    defparam i2022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2023_3_lut (.I0(ram_s_172_7), .I1(sx[7]), .I2(n85), .I3(GND_net), 
            .O(n2271));   // src/ram.vhd(56[12:17])
    defparam i2023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2024_3_lut (.I0(ram_s_173_0), .I1(register_vector[8]), .I2(n84), 
            .I3(GND_net), .O(n2272));   // src/ram.vhd(56[12:17])
    defparam i2024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2025_3_lut (.I0(ram_s_173_1), .I1(register_vector[9]), .I2(n84), 
            .I3(GND_net), .O(n2273));   // src/ram.vhd(56[12:17])
    defparam i2025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2026_3_lut (.I0(ram_s_173_2), .I1(register_vector[10]), .I2(n84), 
            .I3(GND_net), .O(n2274));   // src/ram.vhd(56[12:17])
    defparam i2026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2027_3_lut (.I0(ram_s_173_3), .I1(register_vector[11]), .I2(n84), 
            .I3(GND_net), .O(n2275));   // src/ram.vhd(56[12:17])
    defparam i2027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2028_3_lut (.I0(ram_s_173_4), .I1(sx[4]), .I2(n84), .I3(GND_net), 
            .O(n2276));   // src/ram.vhd(56[12:17])
    defparam i2028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2029_3_lut (.I0(ram_s_173_5), .I1(sx[5]), .I2(n84), .I3(GND_net), 
            .O(n2277));   // src/ram.vhd(56[12:17])
    defparam i2029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2030_3_lut (.I0(ram_s_173_6), .I1(sx[6]), .I2(n84), .I3(GND_net), 
            .O(n2278));   // src/ram.vhd(56[12:17])
    defparam i2030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2031_3_lut (.I0(ram_s_173_7), .I1(sx[7]), .I2(n84), .I3(GND_net), 
            .O(n2279));   // src/ram.vhd(56[12:17])
    defparam i2031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2040_3_lut (.I0(ram_s_175_0), .I1(register_vector[8]), .I2(n82), 
            .I3(GND_net), .O(n2288));   // src/ram.vhd(56[12:17])
    defparam i2040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2041_3_lut (.I0(ram_s_175_1), .I1(register_vector[9]), .I2(n82), 
            .I3(GND_net), .O(n2289));   // src/ram.vhd(56[12:17])
    defparam i2041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2042_3_lut (.I0(ram_s_175_2), .I1(register_vector[10]), .I2(n82), 
            .I3(GND_net), .O(n2290));   // src/ram.vhd(56[12:17])
    defparam i2042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2043_3_lut (.I0(ram_s_175_3), .I1(register_vector[11]), .I2(n82), 
            .I3(GND_net), .O(n2291));   // src/ram.vhd(56[12:17])
    defparam i2043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2044_3_lut (.I0(ram_s_175_4), .I1(sx[4]), .I2(n82), .I3(GND_net), 
            .O(n2292));   // src/ram.vhd(56[12:17])
    defparam i2044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2045_3_lut (.I0(ram_s_175_5), .I1(sx[5]), .I2(n82), .I3(GND_net), 
            .O(n2293));   // src/ram.vhd(56[12:17])
    defparam i2045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2046_3_lut (.I0(ram_s_175_6), .I1(sx[6]), .I2(n82), .I3(GND_net), 
            .O(n2294));   // src/ram.vhd(56[12:17])
    defparam i2046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2047_3_lut (.I0(ram_s_175_7), .I1(sx[7]), .I2(n82), .I3(GND_net), 
            .O(n2295));   // src/ram.vhd(56[12:17])
    defparam i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2120_3_lut (.I0(ram_s_185_0), .I1(register_vector[8]), .I2(n72), 
            .I3(GND_net), .O(n2368));   // src/ram.vhd(56[12:17])
    defparam i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2121_3_lut (.I0(ram_s_185_1), .I1(register_vector[9]), .I2(n72), 
            .I3(GND_net), .O(n2369));   // src/ram.vhd(56[12:17])
    defparam i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2122_3_lut (.I0(ram_s_185_2), .I1(register_vector[10]), .I2(n72), 
            .I3(GND_net), .O(n2370));   // src/ram.vhd(56[12:17])
    defparam i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2123_3_lut (.I0(ram_s_185_3), .I1(register_vector[11]), .I2(n72), 
            .I3(GND_net), .O(n2371));   // src/ram.vhd(56[12:17])
    defparam i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2124_3_lut (.I0(ram_s_185_4), .I1(sx[4]), .I2(n72), .I3(GND_net), 
            .O(n2372));   // src/ram.vhd(56[12:17])
    defparam i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2125_3_lut (.I0(ram_s_185_5), .I1(sx[5]), .I2(n72), .I3(GND_net), 
            .O(n2373));   // src/ram.vhd(56[12:17])
    defparam i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2126_3_lut (.I0(ram_s_185_6), .I1(sx[6]), .I2(n72), .I3(GND_net), 
            .O(n2374));   // src/ram.vhd(56[12:17])
    defparam i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2127_3_lut (.I0(ram_s_185_7), .I1(sx[7]), .I2(n72), .I3(GND_net), 
            .O(n2375));   // src/ram.vhd(56[12:17])
    defparam i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2128_3_lut (.I0(ram_s_186_0), .I1(register_vector[8]), .I2(n71), 
            .I3(GND_net), .O(n2376));   // src/ram.vhd(56[12:17])
    defparam i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2129_3_lut (.I0(ram_s_186_1), .I1(register_vector[9]), .I2(n71), 
            .I3(GND_net), .O(n2377));   // src/ram.vhd(56[12:17])
    defparam i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2130_3_lut (.I0(ram_s_186_2), .I1(register_vector[10]), .I2(n71), 
            .I3(GND_net), .O(n2378));   // src/ram.vhd(56[12:17])
    defparam i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2131_3_lut (.I0(ram_s_186_3), .I1(register_vector[11]), .I2(n71), 
            .I3(GND_net), .O(n2379));   // src/ram.vhd(56[12:17])
    defparam i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2132_3_lut (.I0(ram_s_186_4), .I1(sx[4]), .I2(n71), .I3(GND_net), 
            .O(n2380));   // src/ram.vhd(56[12:17])
    defparam i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2133_3_lut (.I0(ram_s_186_5), .I1(sx[5]), .I2(n71), .I3(GND_net), 
            .O(n2381));   // src/ram.vhd(56[12:17])
    defparam i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2134_3_lut (.I0(ram_s_186_6), .I1(sx[6]), .I2(n71), .I3(GND_net), 
            .O(n2382));   // src/ram.vhd(56[12:17])
    defparam i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2135_3_lut (.I0(ram_s_186_7), .I1(sx[7]), .I2(n71), .I3(GND_net), 
            .O(n2383));   // src/ram.vhd(56[12:17])
    defparam i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2160_3_lut (.I0(ram_s_190_0), .I1(register_vector[8]), .I2(n67), 
            .I3(GND_net), .O(n2408));   // src/ram.vhd(56[12:17])
    defparam i2160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2161_3_lut (.I0(ram_s_190_1), .I1(register_vector[9]), .I2(n67), 
            .I3(GND_net), .O(n2409));   // src/ram.vhd(56[12:17])
    defparam i2161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2162_3_lut (.I0(ram_s_190_2), .I1(register_vector[10]), .I2(n67), 
            .I3(GND_net), .O(n2410));   // src/ram.vhd(56[12:17])
    defparam i2162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2163_3_lut (.I0(ram_s_190_3), .I1(register_vector[11]), .I2(n67), 
            .I3(GND_net), .O(n2411));   // src/ram.vhd(56[12:17])
    defparam i2163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2164_3_lut (.I0(ram_s_190_4), .I1(sx[4]), .I2(n67), .I3(GND_net), 
            .O(n2412));   // src/ram.vhd(56[12:17])
    defparam i2164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2165_3_lut (.I0(ram_s_190_5), .I1(sx[5]), .I2(n67), .I3(GND_net), 
            .O(n2413));   // src/ram.vhd(56[12:17])
    defparam i2165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2166_3_lut (.I0(ram_s_190_6), .I1(sx[6]), .I2(n67), .I3(GND_net), 
            .O(n2414));   // src/ram.vhd(56[12:17])
    defparam i2166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2167_3_lut (.I0(ram_s_190_7), .I1(sx[7]), .I2(n67), .I3(GND_net), 
            .O(n2415));   // src/ram.vhd(56[12:17])
    defparam i2167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2168_3_lut (.I0(ram_s_191_0), .I1(register_vector[8]), .I2(n66), 
            .I3(GND_net), .O(n2416));   // src/ram.vhd(56[12:17])
    defparam i2168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2169_3_lut (.I0(ram_s_191_1), .I1(register_vector[9]), .I2(n66), 
            .I3(GND_net), .O(n2417));   // src/ram.vhd(56[12:17])
    defparam i2169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2170_3_lut (.I0(ram_s_191_2), .I1(register_vector[10]), .I2(n66), 
            .I3(GND_net), .O(n2418));   // src/ram.vhd(56[12:17])
    defparam i2170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2171_3_lut (.I0(ram_s_191_3), .I1(register_vector[11]), .I2(n66), 
            .I3(GND_net), .O(n2419));   // src/ram.vhd(56[12:17])
    defparam i2171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2172_3_lut (.I0(ram_s_191_4), .I1(sx[4]), .I2(n66), .I3(GND_net), 
            .O(n2420));   // src/ram.vhd(56[12:17])
    defparam i2172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2173_3_lut (.I0(ram_s_191_5), .I1(sx[5]), .I2(n66), .I3(GND_net), 
            .O(n2421));   // src/ram.vhd(56[12:17])
    defparam i2173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2174_3_lut (.I0(ram_s_191_6), .I1(sx[6]), .I2(n66), .I3(GND_net), 
            .O(n2422));   // src/ram.vhd(56[12:17])
    defparam i2174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2175_3_lut (.I0(ram_s_191_7), .I1(sx[7]), .I2(n66), .I3(GND_net), 
            .O(n2423));   // src/ram.vhd(56[12:17])
    defparam i2175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2176_3_lut (.I0(ram_s_192_0), .I1(register_vector[8]), .I2(n65), 
            .I3(GND_net), .O(n2424));   // src/ram.vhd(56[12:17])
    defparam i2176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2177_3_lut (.I0(ram_s_192_1), .I1(register_vector[9]), .I2(n65), 
            .I3(GND_net), .O(n2425));   // src/ram.vhd(56[12:17])
    defparam i2177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2178_3_lut (.I0(ram_s_192_2), .I1(register_vector[10]), .I2(n65), 
            .I3(GND_net), .O(n2426));   // src/ram.vhd(56[12:17])
    defparam i2178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2179_3_lut (.I0(ram_s_192_3), .I1(register_vector[11]), .I2(n65), 
            .I3(GND_net), .O(n2427));   // src/ram.vhd(56[12:17])
    defparam i2179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2180_3_lut (.I0(ram_s_192_4), .I1(sx[4]), .I2(n65), .I3(GND_net), 
            .O(n2428));   // src/ram.vhd(56[12:17])
    defparam i2180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2181_3_lut (.I0(ram_s_192_5), .I1(sx[5]), .I2(n65), .I3(GND_net), 
            .O(n2429));   // src/ram.vhd(56[12:17])
    defparam i2181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2182_3_lut (.I0(ram_s_192_6), .I1(sx[6]), .I2(n65), .I3(GND_net), 
            .O(n2430));   // src/ram.vhd(56[12:17])
    defparam i2182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2183_3_lut (.I0(ram_s_192_7), .I1(sx[7]), .I2(n65), .I3(GND_net), 
            .O(n2431));   // src/ram.vhd(56[12:17])
    defparam i2183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2184_3_lut (.I0(ram_s_193_0), .I1(register_vector[8]), .I2(n64), 
            .I3(GND_net), .O(n2432));   // src/ram.vhd(56[12:17])
    defparam i2184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2185_3_lut (.I0(ram_s_193_1), .I1(register_vector[9]), .I2(n64), 
            .I3(GND_net), .O(n2433));   // src/ram.vhd(56[12:17])
    defparam i2185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2186_3_lut (.I0(ram_s_193_2), .I1(register_vector[10]), .I2(n64), 
            .I3(GND_net), .O(n2434));   // src/ram.vhd(56[12:17])
    defparam i2186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2187_3_lut (.I0(ram_s_193_3), .I1(register_vector[11]), .I2(n64), 
            .I3(GND_net), .O(n2435));   // src/ram.vhd(56[12:17])
    defparam i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2188_3_lut (.I0(ram_s_193_4), .I1(sx[4]), .I2(n64), .I3(GND_net), 
            .O(n2436));   // src/ram.vhd(56[12:17])
    defparam i2188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2189_3_lut (.I0(ram_s_193_5), .I1(sx[5]), .I2(n64), .I3(GND_net), 
            .O(n2437));   // src/ram.vhd(56[12:17])
    defparam i2189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2190_3_lut (.I0(ram_s_193_6), .I1(sx[6]), .I2(n64), .I3(GND_net), 
            .O(n2438));   // src/ram.vhd(56[12:17])
    defparam i2190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2191_3_lut (.I0(ram_s_193_7), .I1(sx[7]), .I2(n64), .I3(GND_net), 
            .O(n2439));   // src/ram.vhd(56[12:17])
    defparam i2191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2192_3_lut (.I0(ram_s_194_0), .I1(register_vector[8]), .I2(n63), 
            .I3(GND_net), .O(n2440));   // src/ram.vhd(56[12:17])
    defparam i2192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2193_3_lut (.I0(ram_s_194_1), .I1(register_vector[9]), .I2(n63), 
            .I3(GND_net), .O(n2441));   // src/ram.vhd(56[12:17])
    defparam i2193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2194_3_lut (.I0(ram_s_194_2), .I1(register_vector[10]), .I2(n63), 
            .I3(GND_net), .O(n2442));   // src/ram.vhd(56[12:17])
    defparam i2194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2195_3_lut (.I0(ram_s_194_3), .I1(register_vector[11]), .I2(n63), 
            .I3(GND_net), .O(n2443));   // src/ram.vhd(56[12:17])
    defparam i2195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2196_3_lut (.I0(ram_s_194_4), .I1(sx[4]), .I2(n63), .I3(GND_net), 
            .O(n2444));   // src/ram.vhd(56[12:17])
    defparam i2196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2197_3_lut (.I0(ram_s_194_5), .I1(sx[5]), .I2(n63), .I3(GND_net), 
            .O(n2445));   // src/ram.vhd(56[12:17])
    defparam i2197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2198_3_lut (.I0(ram_s_194_6), .I1(sx[6]), .I2(n63), .I3(GND_net), 
            .O(n2446));   // src/ram.vhd(56[12:17])
    defparam i2198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2199_3_lut (.I0(ram_s_194_7), .I1(sx[7]), .I2(n63), .I3(GND_net), 
            .O(n2447));   // src/ram.vhd(56[12:17])
    defparam i2199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2200_3_lut (.I0(ram_s_195_0), .I1(register_vector[8]), .I2(n62), 
            .I3(GND_net), .O(n2448));   // src/ram.vhd(56[12:17])
    defparam i2200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2201_3_lut (.I0(ram_s_195_1), .I1(register_vector[9]), .I2(n62), 
            .I3(GND_net), .O(n2449));   // src/ram.vhd(56[12:17])
    defparam i2201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2202_3_lut (.I0(ram_s_195_2), .I1(register_vector[10]), .I2(n62), 
            .I3(GND_net), .O(n2450));   // src/ram.vhd(56[12:17])
    defparam i2202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2203_3_lut (.I0(ram_s_195_3), .I1(register_vector[11]), .I2(n62), 
            .I3(GND_net), .O(n2451));   // src/ram.vhd(56[12:17])
    defparam i2203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2204_3_lut (.I0(ram_s_195_4), .I1(sx[4]), .I2(n62), .I3(GND_net), 
            .O(n2452));   // src/ram.vhd(56[12:17])
    defparam i2204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2205_3_lut (.I0(ram_s_195_5), .I1(sx[5]), .I2(n62), .I3(GND_net), 
            .O(n2453));   // src/ram.vhd(56[12:17])
    defparam i2205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2206_3_lut (.I0(ram_s_195_6), .I1(sx[6]), .I2(n62), .I3(GND_net), 
            .O(n2454));   // src/ram.vhd(56[12:17])
    defparam i2206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2207_3_lut (.I0(ram_s_195_7), .I1(sx[7]), .I2(n62), .I3(GND_net), 
            .O(n2455));   // src/ram.vhd(56[12:17])
    defparam i2207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2208_3_lut (.I0(ram_s_196_0), .I1(register_vector[8]), .I2(n61), 
            .I3(GND_net), .O(n2456));   // src/ram.vhd(56[12:17])
    defparam i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2209_3_lut (.I0(ram_s_196_1), .I1(register_vector[9]), .I2(n61), 
            .I3(GND_net), .O(n2457));   // src/ram.vhd(56[12:17])
    defparam i2209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2210_3_lut (.I0(ram_s_196_2), .I1(register_vector[10]), .I2(n61), 
            .I3(GND_net), .O(n2458));   // src/ram.vhd(56[12:17])
    defparam i2210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2211_3_lut (.I0(ram_s_196_3), .I1(register_vector[11]), .I2(n61), 
            .I3(GND_net), .O(n2459));   // src/ram.vhd(56[12:17])
    defparam i2211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2212_3_lut (.I0(ram_s_196_4), .I1(sx[4]), .I2(n61), .I3(GND_net), 
            .O(n2460));   // src/ram.vhd(56[12:17])
    defparam i2212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2213_3_lut (.I0(ram_s_196_5), .I1(sx[5]), .I2(n61), .I3(GND_net), 
            .O(n2461));   // src/ram.vhd(56[12:17])
    defparam i2213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2214_3_lut (.I0(ram_s_196_6), .I1(sx[6]), .I2(n61), .I3(GND_net), 
            .O(n2462));   // src/ram.vhd(56[12:17])
    defparam i2214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2215_3_lut (.I0(ram_s_196_7), .I1(sx[7]), .I2(n61), .I3(GND_net), 
            .O(n2463));   // src/ram.vhd(56[12:17])
    defparam i2215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2216_3_lut (.I0(ram_s_197_0), .I1(register_vector[8]), .I2(n60), 
            .I3(GND_net), .O(n2464));   // src/ram.vhd(56[12:17])
    defparam i2216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2217_3_lut (.I0(ram_s_197_1), .I1(register_vector[9]), .I2(n60), 
            .I3(GND_net), .O(n2465));   // src/ram.vhd(56[12:17])
    defparam i2217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2218_3_lut (.I0(ram_s_197_2), .I1(register_vector[10]), .I2(n60), 
            .I3(GND_net), .O(n2466));   // src/ram.vhd(56[12:17])
    defparam i2218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2219_3_lut (.I0(ram_s_197_3), .I1(register_vector[11]), .I2(n60), 
            .I3(GND_net), .O(n2467));   // src/ram.vhd(56[12:17])
    defparam i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2220_3_lut (.I0(ram_s_197_4), .I1(sx[4]), .I2(n60), .I3(GND_net), 
            .O(n2468));   // src/ram.vhd(56[12:17])
    defparam i2220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2221_3_lut (.I0(ram_s_197_5), .I1(sx[5]), .I2(n60), .I3(GND_net), 
            .O(n2469));   // src/ram.vhd(56[12:17])
    defparam i2221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2222_3_lut (.I0(ram_s_197_6), .I1(sx[6]), .I2(n60), .I3(GND_net), 
            .O(n2470));   // src/ram.vhd(56[12:17])
    defparam i2222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2223_3_lut (.I0(ram_s_197_7), .I1(sx[7]), .I2(n60), .I3(GND_net), 
            .O(n2471));   // src/ram.vhd(56[12:17])
    defparam i2223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2224_3_lut (.I0(ram_s_198_0), .I1(register_vector[8]), .I2(n59), 
            .I3(GND_net), .O(n2472));   // src/ram.vhd(56[12:17])
    defparam i2224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2225_3_lut (.I0(ram_s_198_1), .I1(register_vector[9]), .I2(n59), 
            .I3(GND_net), .O(n2473));   // src/ram.vhd(56[12:17])
    defparam i2225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2226_3_lut (.I0(ram_s_198_2), .I1(register_vector[10]), .I2(n59), 
            .I3(GND_net), .O(n2474));   // src/ram.vhd(56[12:17])
    defparam i2226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2227_3_lut (.I0(ram_s_198_3), .I1(register_vector[11]), .I2(n59), 
            .I3(GND_net), .O(n2475));   // src/ram.vhd(56[12:17])
    defparam i2227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2228_3_lut (.I0(ram_s_198_4), .I1(sx[4]), .I2(n59), .I3(GND_net), 
            .O(n2476));   // src/ram.vhd(56[12:17])
    defparam i2228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2229_3_lut (.I0(ram_s_198_5), .I1(sx[5]), .I2(n59), .I3(GND_net), 
            .O(n2477));   // src/ram.vhd(56[12:17])
    defparam i2229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2230_3_lut (.I0(ram_s_198_6), .I1(sx[6]), .I2(n59), .I3(GND_net), 
            .O(n2478));   // src/ram.vhd(56[12:17])
    defparam i2230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2231_3_lut (.I0(ram_s_198_7), .I1(sx[7]), .I2(n59), .I3(GND_net), 
            .O(n2479));   // src/ram.vhd(56[12:17])
    defparam i2231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2232_3_lut (.I0(ram_s_199_0), .I1(register_vector[8]), .I2(n58), 
            .I3(GND_net), .O(n2480));   // src/ram.vhd(56[12:17])
    defparam i2232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2233_3_lut (.I0(ram_s_199_1), .I1(register_vector[9]), .I2(n58), 
            .I3(GND_net), .O(n2481));   // src/ram.vhd(56[12:17])
    defparam i2233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2234_3_lut (.I0(ram_s_199_2), .I1(register_vector[10]), .I2(n58), 
            .I3(GND_net), .O(n2482));   // src/ram.vhd(56[12:17])
    defparam i2234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2235_3_lut (.I0(ram_s_199_3), .I1(register_vector[11]), .I2(n58), 
            .I3(GND_net), .O(n2483));   // src/ram.vhd(56[12:17])
    defparam i2235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2236_3_lut (.I0(ram_s_199_4), .I1(sx[4]), .I2(n58), .I3(GND_net), 
            .O(n2484));   // src/ram.vhd(56[12:17])
    defparam i2236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2237_3_lut (.I0(ram_s_199_5), .I1(sx[5]), .I2(n58), .I3(GND_net), 
            .O(n2485));   // src/ram.vhd(56[12:17])
    defparam i2237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2238_3_lut (.I0(ram_s_199_6), .I1(sx[6]), .I2(n58), .I3(GND_net), 
            .O(n2486));   // src/ram.vhd(56[12:17])
    defparam i2238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2239_3_lut (.I0(ram_s_199_7), .I1(sx[7]), .I2(n58), .I3(GND_net), 
            .O(n2487));   // src/ram.vhd(56[12:17])
    defparam i2239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2240_3_lut (.I0(ram_s_200_0), .I1(register_vector[8]), .I2(n57), 
            .I3(GND_net), .O(n2488));   // src/ram.vhd(56[12:17])
    defparam i2240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2241_3_lut (.I0(ram_s_200_1), .I1(register_vector[9]), .I2(n57), 
            .I3(GND_net), .O(n2489));   // src/ram.vhd(56[12:17])
    defparam i2241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2242_3_lut (.I0(ram_s_200_2), .I1(register_vector[10]), .I2(n57), 
            .I3(GND_net), .O(n2490));   // src/ram.vhd(56[12:17])
    defparam i2242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2243_3_lut (.I0(ram_s_200_3), .I1(register_vector[11]), .I2(n57), 
            .I3(GND_net), .O(n2491));   // src/ram.vhd(56[12:17])
    defparam i2243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2244_3_lut (.I0(ram_s_200_4), .I1(sx[4]), .I2(n57), .I3(GND_net), 
            .O(n2492));   // src/ram.vhd(56[12:17])
    defparam i2244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2245_3_lut (.I0(ram_s_200_5), .I1(sx[5]), .I2(n57), .I3(GND_net), 
            .O(n2493));   // src/ram.vhd(56[12:17])
    defparam i2245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2246_3_lut (.I0(ram_s_200_6), .I1(sx[6]), .I2(n57), .I3(GND_net), 
            .O(n2494));   // src/ram.vhd(56[12:17])
    defparam i2246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2247_3_lut (.I0(ram_s_200_7), .I1(sx[7]), .I2(n57), .I3(GND_net), 
            .O(n2495));   // src/ram.vhd(56[12:17])
    defparam i2247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2248_3_lut (.I0(ram_s_201_0), .I1(register_vector[8]), .I2(n56), 
            .I3(GND_net), .O(n2496));   // src/ram.vhd(56[12:17])
    defparam i2248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2249_3_lut (.I0(ram_s_201_1), .I1(register_vector[9]), .I2(n56), 
            .I3(GND_net), .O(n2497));   // src/ram.vhd(56[12:17])
    defparam i2249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2250_3_lut (.I0(ram_s_201_2), .I1(register_vector[10]), .I2(n56), 
            .I3(GND_net), .O(n2498));   // src/ram.vhd(56[12:17])
    defparam i2250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2251_3_lut (.I0(ram_s_201_3), .I1(register_vector[11]), .I2(n56), 
            .I3(GND_net), .O(n2499));   // src/ram.vhd(56[12:17])
    defparam i2251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2252_3_lut (.I0(ram_s_201_4), .I1(sx[4]), .I2(n56), .I3(GND_net), 
            .O(n2500));   // src/ram.vhd(56[12:17])
    defparam i2252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2253_3_lut (.I0(ram_s_201_5), .I1(sx[5]), .I2(n56), .I3(GND_net), 
            .O(n2501));   // src/ram.vhd(56[12:17])
    defparam i2253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2254_3_lut (.I0(ram_s_201_6), .I1(sx[6]), .I2(n56), .I3(GND_net), 
            .O(n2502));   // src/ram.vhd(56[12:17])
    defparam i2254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2255_3_lut (.I0(ram_s_201_7), .I1(sx[7]), .I2(n56), .I3(GND_net), 
            .O(n2503));   // src/ram.vhd(56[12:17])
    defparam i2255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2256_3_lut (.I0(ram_s_202_0), .I1(register_vector[8]), .I2(n55), 
            .I3(GND_net), .O(n2504));   // src/ram.vhd(56[12:17])
    defparam i2256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2257_3_lut (.I0(ram_s_202_1), .I1(register_vector[9]), .I2(n55), 
            .I3(GND_net), .O(n2505));   // src/ram.vhd(56[12:17])
    defparam i2257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2258_3_lut (.I0(ram_s_202_2), .I1(register_vector[10]), .I2(n55), 
            .I3(GND_net), .O(n2506));   // src/ram.vhd(56[12:17])
    defparam i2258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2259_3_lut (.I0(ram_s_202_3), .I1(register_vector[11]), .I2(n55), 
            .I3(GND_net), .O(n2507));   // src/ram.vhd(56[12:17])
    defparam i2259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2260_3_lut (.I0(ram_s_202_4), .I1(sx[4]), .I2(n55), .I3(GND_net), 
            .O(n2508));   // src/ram.vhd(56[12:17])
    defparam i2260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2261_3_lut (.I0(ram_s_202_5), .I1(sx[5]), .I2(n55), .I3(GND_net), 
            .O(n2509));   // src/ram.vhd(56[12:17])
    defparam i2261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2262_3_lut (.I0(ram_s_202_6), .I1(sx[6]), .I2(n55), .I3(GND_net), 
            .O(n2510));   // src/ram.vhd(56[12:17])
    defparam i2262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2263_3_lut (.I0(ram_s_202_7), .I1(sx[7]), .I2(n55), .I3(GND_net), 
            .O(n2511));   // src/ram.vhd(56[12:17])
    defparam i2263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2264_3_lut (.I0(ram_s_203_0), .I1(register_vector[8]), .I2(n54), 
            .I3(GND_net), .O(n2512));   // src/ram.vhd(56[12:17])
    defparam i2264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2265_3_lut (.I0(ram_s_203_1), .I1(register_vector[9]), .I2(n54), 
            .I3(GND_net), .O(n2513));   // src/ram.vhd(56[12:17])
    defparam i2265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2266_3_lut (.I0(ram_s_203_2), .I1(register_vector[10]), .I2(n54), 
            .I3(GND_net), .O(n2514));   // src/ram.vhd(56[12:17])
    defparam i2266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2267_3_lut (.I0(ram_s_203_3), .I1(register_vector[11]), .I2(n54), 
            .I3(GND_net), .O(n2515));   // src/ram.vhd(56[12:17])
    defparam i2267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2268_3_lut (.I0(ram_s_203_4), .I1(sx[4]), .I2(n54), .I3(GND_net), 
            .O(n2516));   // src/ram.vhd(56[12:17])
    defparam i2268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2269_3_lut (.I0(ram_s_203_5), .I1(sx[5]), .I2(n54), .I3(GND_net), 
            .O(n2517));   // src/ram.vhd(56[12:17])
    defparam i2269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2270_3_lut (.I0(ram_s_203_6), .I1(sx[6]), .I2(n54), .I3(GND_net), 
            .O(n2518));   // src/ram.vhd(56[12:17])
    defparam i2270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2271_3_lut (.I0(ram_s_203_7), .I1(sx[7]), .I2(n54), .I3(GND_net), 
            .O(n2519));   // src/ram.vhd(56[12:17])
    defparam i2271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1247_3_lut (.I0(ram_s_75_7), .I1(sx[7]), .I2(n182), .I3(GND_net), 
            .O(n1495));   // src/ram.vhd(56[12:17])
    defparam i1247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1246_3_lut (.I0(ram_s_75_6), .I1(sx[6]), .I2(n182), .I3(GND_net), 
            .O(n1494));   // src/ram.vhd(56[12:17])
    defparam i1246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1245_3_lut (.I0(ram_s_75_5), .I1(sx[5]), .I2(n182), .I3(GND_net), 
            .O(n1493));   // src/ram.vhd(56[12:17])
    defparam i1245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1244_3_lut (.I0(ram_s_75_4), .I1(sx[4]), .I2(n182), .I3(GND_net), 
            .O(n1492));   // src/ram.vhd(56[12:17])
    defparam i1244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1243_3_lut (.I0(ram_s_75_3), .I1(register_vector[11]), .I2(n182), 
            .I3(GND_net), .O(n1491));   // src/ram.vhd(56[12:17])
    defparam i1243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1242_3_lut (.I0(ram_s_75_2), .I1(register_vector[10]), .I2(n182), 
            .I3(GND_net), .O(n1490));   // src/ram.vhd(56[12:17])
    defparam i1242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1241_3_lut (.I0(ram_s_75_1), .I1(register_vector[9]), .I2(n182), 
            .I3(GND_net), .O(n1489));   // src/ram.vhd(56[12:17])
    defparam i1241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1240_3_lut (.I0(ram_s_75_0), .I1(register_vector[8]), .I2(n182), 
            .I3(GND_net), .O(n1488));   // src/ram.vhd(56[12:17])
    defparam i1240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1239_3_lut (.I0(ram_s_74_7), .I1(sx[7]), .I2(n183), .I3(GND_net), 
            .O(n1487));   // src/ram.vhd(56[12:17])
    defparam i1239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1238_3_lut (.I0(ram_s_74_6), .I1(sx[6]), .I2(n183), .I3(GND_net), 
            .O(n1486));   // src/ram.vhd(56[12:17])
    defparam i1238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1237_3_lut (.I0(ram_s_74_5), .I1(sx[5]), .I2(n183), .I3(GND_net), 
            .O(n1485));   // src/ram.vhd(56[12:17])
    defparam i1237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1236_3_lut (.I0(ram_s_74_4), .I1(sx[4]), .I2(n183), .I3(GND_net), 
            .O(n1484));   // src/ram.vhd(56[12:17])
    defparam i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1235_3_lut (.I0(ram_s_74_3), .I1(register_vector[11]), .I2(n183), 
            .I3(GND_net), .O(n1483));   // src/ram.vhd(56[12:17])
    defparam i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1234_3_lut (.I0(ram_s_74_2), .I1(register_vector[10]), .I2(n183), 
            .I3(GND_net), .O(n1482));   // src/ram.vhd(56[12:17])
    defparam i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1233_3_lut (.I0(ram_s_74_1), .I1(register_vector[9]), .I2(n183), 
            .I3(GND_net), .O(n1481));   // src/ram.vhd(56[12:17])
    defparam i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1232_3_lut (.I0(ram_s_74_0), .I1(register_vector[8]), .I2(n183), 
            .I3(GND_net), .O(n1480));   // src/ram.vhd(56[12:17])
    defparam i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1231_3_lut (.I0(ram_s_73_7), .I1(sx[7]), .I2(n184), .I3(GND_net), 
            .O(n1479));   // src/ram.vhd(56[12:17])
    defparam i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1230_3_lut (.I0(ram_s_73_6), .I1(sx[6]), .I2(n184), .I3(GND_net), 
            .O(n1478));   // src/ram.vhd(56[12:17])
    defparam i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1229_3_lut (.I0(ram_s_73_5), .I1(sx[5]), .I2(n184), .I3(GND_net), 
            .O(n1477));   // src/ram.vhd(56[12:17])
    defparam i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1228_3_lut (.I0(ram_s_73_4), .I1(sx[4]), .I2(n184), .I3(GND_net), 
            .O(n1476));   // src/ram.vhd(56[12:17])
    defparam i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1227_3_lut (.I0(ram_s_73_3), .I1(register_vector[11]), .I2(n184), 
            .I3(GND_net), .O(n1475));   // src/ram.vhd(56[12:17])
    defparam i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1226_3_lut (.I0(ram_s_73_2), .I1(register_vector[10]), .I2(n184), 
            .I3(GND_net), .O(n1474));   // src/ram.vhd(56[12:17])
    defparam i1226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1225_3_lut (.I0(ram_s_73_1), .I1(register_vector[9]), .I2(n184), 
            .I3(GND_net), .O(n1473));   // src/ram.vhd(56[12:17])
    defparam i1225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1224_3_lut (.I0(ram_s_73_0), .I1(register_vector[8]), .I2(n184), 
            .I3(GND_net), .O(n1472));   // src/ram.vhd(56[12:17])
    defparam i1224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1223_3_lut (.I0(ram_s_72_7), .I1(sx[7]), .I2(n185), .I3(GND_net), 
            .O(n1471));   // src/ram.vhd(56[12:17])
    defparam i1223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1222_3_lut (.I0(ram_s_72_6), .I1(sx[6]), .I2(n185), .I3(GND_net), 
            .O(n1470));   // src/ram.vhd(56[12:17])
    defparam i1222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1221_3_lut (.I0(ram_s_72_5), .I1(sx[5]), .I2(n185), .I3(GND_net), 
            .O(n1469));   // src/ram.vhd(56[12:17])
    defparam i1221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1220_3_lut (.I0(ram_s_72_4), .I1(sx[4]), .I2(n185), .I3(GND_net), 
            .O(n1468));   // src/ram.vhd(56[12:17])
    defparam i1220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1219_3_lut (.I0(ram_s_72_3), .I1(register_vector[11]), .I2(n185), 
            .I3(GND_net), .O(n1467));   // src/ram.vhd(56[12:17])
    defparam i1219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1218_3_lut (.I0(ram_s_72_2), .I1(register_vector[10]), .I2(n185), 
            .I3(GND_net), .O(n1466));   // src/ram.vhd(56[12:17])
    defparam i1218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1217_3_lut (.I0(ram_s_72_1), .I1(register_vector[9]), .I2(n185), 
            .I3(GND_net), .O(n1465));   // src/ram.vhd(56[12:17])
    defparam i1217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1216_3_lut (.I0(ram_s_72_0), .I1(register_vector[8]), .I2(n185), 
            .I3(GND_net), .O(n1464));   // src/ram.vhd(56[12:17])
    defparam i1216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1215_3_lut (.I0(ram_s_71_7), .I1(sx[7]), .I2(n186), .I3(GND_net), 
            .O(n1463));   // src/ram.vhd(56[12:17])
    defparam i1215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1214_3_lut (.I0(ram_s_71_6), .I1(sx[6]), .I2(n186), .I3(GND_net), 
            .O(n1462));   // src/ram.vhd(56[12:17])
    defparam i1214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1213_3_lut (.I0(ram_s_71_5), .I1(sx[5]), .I2(n186), .I3(GND_net), 
            .O(n1461));   // src/ram.vhd(56[12:17])
    defparam i1213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1212_3_lut (.I0(ram_s_71_4), .I1(sx[4]), .I2(n186), .I3(GND_net), 
            .O(n1460));   // src/ram.vhd(56[12:17])
    defparam i1212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1211_3_lut (.I0(ram_s_71_3), .I1(register_vector[11]), .I2(n186), 
            .I3(GND_net), .O(n1459));   // src/ram.vhd(56[12:17])
    defparam i1211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1210_3_lut (.I0(ram_s_71_2), .I1(register_vector[10]), .I2(n186), 
            .I3(GND_net), .O(n1458));   // src/ram.vhd(56[12:17])
    defparam i1210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1209_3_lut (.I0(ram_s_71_1), .I1(register_vector[9]), .I2(n186), 
            .I3(GND_net), .O(n1457));   // src/ram.vhd(56[12:17])
    defparam i1209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1208_3_lut (.I0(ram_s_71_0), .I1(register_vector[8]), .I2(n186), 
            .I3(GND_net), .O(n1456));   // src/ram.vhd(56[12:17])
    defparam i1208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1207_3_lut (.I0(ram_s_70_7), .I1(sx[7]), .I2(n187), .I3(GND_net), 
            .O(n1455));   // src/ram.vhd(56[12:17])
    defparam i1207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1206_3_lut (.I0(ram_s_70_6), .I1(sx[6]), .I2(n187), .I3(GND_net), 
            .O(n1454));   // src/ram.vhd(56[12:17])
    defparam i1206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1205_3_lut (.I0(ram_s_70_5), .I1(sx[5]), .I2(n187), .I3(GND_net), 
            .O(n1453));   // src/ram.vhd(56[12:17])
    defparam i1205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1204_3_lut (.I0(ram_s_70_4), .I1(sx[4]), .I2(n187), .I3(GND_net), 
            .O(n1452));   // src/ram.vhd(56[12:17])
    defparam i1204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1203_3_lut (.I0(ram_s_70_3), .I1(register_vector[11]), .I2(n187), 
            .I3(GND_net), .O(n1451));   // src/ram.vhd(56[12:17])
    defparam i1203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1202_3_lut (.I0(ram_s_70_2), .I1(register_vector[10]), .I2(n187), 
            .I3(GND_net), .O(n1450));   // src/ram.vhd(56[12:17])
    defparam i1202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1201_3_lut (.I0(ram_s_70_1), .I1(register_vector[9]), .I2(n187), 
            .I3(GND_net), .O(n1449));   // src/ram.vhd(56[12:17])
    defparam i1201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1200_3_lut (.I0(ram_s_70_0), .I1(register_vector[8]), .I2(n187), 
            .I3(GND_net), .O(n1448));   // src/ram.vhd(56[12:17])
    defparam i1200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1199_3_lut (.I0(ram_s_69_7), .I1(sx[7]), .I2(n188), .I3(GND_net), 
            .O(n1447));   // src/ram.vhd(56[12:17])
    defparam i1199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1198_3_lut (.I0(ram_s_69_6), .I1(sx[6]), .I2(n188), .I3(GND_net), 
            .O(n1446));   // src/ram.vhd(56[12:17])
    defparam i1198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1197_3_lut (.I0(ram_s_69_5), .I1(sx[5]), .I2(n188), .I3(GND_net), 
            .O(n1445));   // src/ram.vhd(56[12:17])
    defparam i1197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1196_3_lut (.I0(ram_s_69_4), .I1(sx[4]), .I2(n188), .I3(GND_net), 
            .O(n1444));   // src/ram.vhd(56[12:17])
    defparam i1196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1195_3_lut (.I0(ram_s_69_3), .I1(register_vector[11]), .I2(n188), 
            .I3(GND_net), .O(n1443));   // src/ram.vhd(56[12:17])
    defparam i1195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1194_3_lut (.I0(ram_s_69_2), .I1(register_vector[10]), .I2(n188), 
            .I3(GND_net), .O(n1442));   // src/ram.vhd(56[12:17])
    defparam i1194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1193_3_lut (.I0(ram_s_69_1), .I1(register_vector[9]), .I2(n188), 
            .I3(GND_net), .O(n1441));   // src/ram.vhd(56[12:17])
    defparam i1193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1192_3_lut (.I0(ram_s_69_0), .I1(register_vector[8]), .I2(n188), 
            .I3(GND_net), .O(n1440));   // src/ram.vhd(56[12:17])
    defparam i1192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1191_3_lut (.I0(ram_s_68_7), .I1(sx[7]), .I2(n189), .I3(GND_net), 
            .O(n1439));   // src/ram.vhd(56[12:17])
    defparam i1191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1190_3_lut (.I0(ram_s_68_6), .I1(sx[6]), .I2(n189), .I3(GND_net), 
            .O(n1438));   // src/ram.vhd(56[12:17])
    defparam i1190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1189_3_lut (.I0(ram_s_68_5), .I1(sx[5]), .I2(n189), .I3(GND_net), 
            .O(n1437));   // src/ram.vhd(56[12:17])
    defparam i1189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1188_3_lut (.I0(ram_s_68_4), .I1(sx[4]), .I2(n189), .I3(GND_net), 
            .O(n1436));   // src/ram.vhd(56[12:17])
    defparam i1188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1187_3_lut (.I0(ram_s_68_3), .I1(register_vector[11]), .I2(n189), 
            .I3(GND_net), .O(n1435));   // src/ram.vhd(56[12:17])
    defparam i1187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1186_3_lut (.I0(ram_s_68_2), .I1(register_vector[10]), .I2(n189), 
            .I3(GND_net), .O(n1434));   // src/ram.vhd(56[12:17])
    defparam i1186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1185_3_lut (.I0(ram_s_68_1), .I1(register_vector[9]), .I2(n189), 
            .I3(GND_net), .O(n1433));   // src/ram.vhd(56[12:17])
    defparam i1185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1184_3_lut (.I0(ram_s_68_0), .I1(register_vector[8]), .I2(n189), 
            .I3(GND_net), .O(n1432));   // src/ram.vhd(56[12:17])
    defparam i1184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1183_3_lut (.I0(ram_s_67_7), .I1(sx[7]), .I2(n190), .I3(GND_net), 
            .O(n1431));   // src/ram.vhd(56[12:17])
    defparam i1183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1182_3_lut (.I0(ram_s_67_6), .I1(sx[6]), .I2(n190), .I3(GND_net), 
            .O(n1430));   // src/ram.vhd(56[12:17])
    defparam i1182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1181_3_lut (.I0(ram_s_67_5), .I1(sx[5]), .I2(n190), .I3(GND_net), 
            .O(n1429));   // src/ram.vhd(56[12:17])
    defparam i1181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1180_3_lut (.I0(ram_s_67_4), .I1(sx[4]), .I2(n190), .I3(GND_net), 
            .O(n1428));   // src/ram.vhd(56[12:17])
    defparam i1180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1179_3_lut (.I0(ram_s_67_3), .I1(register_vector[11]), .I2(n190), 
            .I3(GND_net), .O(n1427));   // src/ram.vhd(56[12:17])
    defparam i1179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1178_3_lut (.I0(ram_s_67_2), .I1(register_vector[10]), .I2(n190), 
            .I3(GND_net), .O(n1426));   // src/ram.vhd(56[12:17])
    defparam i1178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1177_3_lut (.I0(ram_s_67_1), .I1(register_vector[9]), .I2(n190), 
            .I3(GND_net), .O(n1425));   // src/ram.vhd(56[12:17])
    defparam i1177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1176_3_lut (.I0(ram_s_67_0), .I1(register_vector[8]), .I2(n190), 
            .I3(GND_net), .O(n1424));   // src/ram.vhd(56[12:17])
    defparam i1176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1175_3_lut (.I0(ram_s_66_7), .I1(sx[7]), .I2(n191), .I3(GND_net), 
            .O(n1423));   // src/ram.vhd(56[12:17])
    defparam i1175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1174_3_lut (.I0(ram_s_66_6), .I1(sx[6]), .I2(n191), .I3(GND_net), 
            .O(n1422));   // src/ram.vhd(56[12:17])
    defparam i1174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1173_3_lut (.I0(ram_s_66_5), .I1(sx[5]), .I2(n191), .I3(GND_net), 
            .O(n1421));   // src/ram.vhd(56[12:17])
    defparam i1173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1172_3_lut (.I0(ram_s_66_4), .I1(sx[4]), .I2(n191), .I3(GND_net), 
            .O(n1420));   // src/ram.vhd(56[12:17])
    defparam i1172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1171_3_lut (.I0(ram_s_66_3), .I1(register_vector[11]), .I2(n191), 
            .I3(GND_net), .O(n1419));   // src/ram.vhd(56[12:17])
    defparam i1171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1170_3_lut (.I0(ram_s_66_2), .I1(register_vector[10]), .I2(n191), 
            .I3(GND_net), .O(n1418));   // src/ram.vhd(56[12:17])
    defparam i1170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1169_3_lut (.I0(ram_s_66_1), .I1(register_vector[9]), .I2(n191), 
            .I3(GND_net), .O(n1417));   // src/ram.vhd(56[12:17])
    defparam i1169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1168_3_lut (.I0(ram_s_66_0), .I1(register_vector[8]), .I2(n191), 
            .I3(GND_net), .O(n1416));   // src/ram.vhd(56[12:17])
    defparam i1168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1167_3_lut (.I0(ram_s_65_7), .I1(sx[7]), .I2(n192), .I3(GND_net), 
            .O(n1415));   // src/ram.vhd(56[12:17])
    defparam i1167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1166_3_lut (.I0(ram_s_65_6), .I1(sx[6]), .I2(n192), .I3(GND_net), 
            .O(n1414));   // src/ram.vhd(56[12:17])
    defparam i1166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1165_3_lut (.I0(ram_s_65_5), .I1(sx[5]), .I2(n192), .I3(GND_net), 
            .O(n1413));   // src/ram.vhd(56[12:17])
    defparam i1165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1164_3_lut (.I0(ram_s_65_4), .I1(sx[4]), .I2(n192), .I3(GND_net), 
            .O(n1412));   // src/ram.vhd(56[12:17])
    defparam i1164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1163_3_lut (.I0(ram_s_65_3), .I1(register_vector[11]), .I2(n192), 
            .I3(GND_net), .O(n1411));   // src/ram.vhd(56[12:17])
    defparam i1163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1162_3_lut (.I0(ram_s_65_2), .I1(register_vector[10]), .I2(n192), 
            .I3(GND_net), .O(n1410));   // src/ram.vhd(56[12:17])
    defparam i1162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1161_3_lut (.I0(ram_s_65_1), .I1(register_vector[9]), .I2(n192), 
            .I3(GND_net), .O(n1409));   // src/ram.vhd(56[12:17])
    defparam i1161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1160_3_lut (.I0(ram_s_65_0), .I1(register_vector[8]), .I2(n192), 
            .I3(GND_net), .O(n1408));   // src/ram.vhd(56[12:17])
    defparam i1160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1159_3_lut (.I0(ram_s_64_7), .I1(sx[7]), .I2(n193), .I3(GND_net), 
            .O(n1407));   // src/ram.vhd(56[12:17])
    defparam i1159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1158_3_lut (.I0(ram_s_64_6), .I1(sx[6]), .I2(n193), .I3(GND_net), 
            .O(n1406));   // src/ram.vhd(56[12:17])
    defparam i1158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1157_3_lut (.I0(ram_s_64_5), .I1(sx[5]), .I2(n193), .I3(GND_net), 
            .O(n1405));   // src/ram.vhd(56[12:17])
    defparam i1157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1156_3_lut (.I0(ram_s_64_4), .I1(sx[4]), .I2(n193), .I3(GND_net), 
            .O(n1404));   // src/ram.vhd(56[12:17])
    defparam i1156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1155_3_lut (.I0(ram_s_64_3), .I1(register_vector[11]), .I2(n193), 
            .I3(GND_net), .O(n1403));   // src/ram.vhd(56[12:17])
    defparam i1155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1154_3_lut (.I0(ram_s_64_2), .I1(register_vector[10]), .I2(n193), 
            .I3(GND_net), .O(n1402));   // src/ram.vhd(56[12:17])
    defparam i1154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1153_3_lut (.I0(ram_s_64_1), .I1(register_vector[9]), .I2(n193), 
            .I3(GND_net), .O(n1401));   // src/ram.vhd(56[12:17])
    defparam i1153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1152_3_lut (.I0(ram_s_64_0), .I1(register_vector[8]), .I2(n193), 
            .I3(GND_net), .O(n1400));   // src/ram.vhd(56[12:17])
    defparam i1152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1151_3_lut (.I0(ram_s_63_7), .I1(sx[7]), .I2(n194), .I3(GND_net), 
            .O(n1399));   // src/ram.vhd(56[12:17])
    defparam i1151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1150_3_lut (.I0(ram_s_63_6), .I1(sx[6]), .I2(n194), .I3(GND_net), 
            .O(n1398));   // src/ram.vhd(56[12:17])
    defparam i1150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1149_3_lut (.I0(ram_s_63_5), .I1(sx[5]), .I2(n194), .I3(GND_net), 
            .O(n1397));   // src/ram.vhd(56[12:17])
    defparam i1149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1148_3_lut (.I0(ram_s_63_4), .I1(sx[4]), .I2(n194), .I3(GND_net), 
            .O(n1396));   // src/ram.vhd(56[12:17])
    defparam i1148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1147_3_lut (.I0(ram_s_63_3), .I1(register_vector[11]), .I2(n194), 
            .I3(GND_net), .O(n1395));   // src/ram.vhd(56[12:17])
    defparam i1147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1146_3_lut (.I0(ram_s_63_2), .I1(register_vector[10]), .I2(n194), 
            .I3(GND_net), .O(n1394));   // src/ram.vhd(56[12:17])
    defparam i1146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1145_3_lut (.I0(ram_s_63_1), .I1(register_vector[9]), .I2(n194), 
            .I3(GND_net), .O(n1393));   // src/ram.vhd(56[12:17])
    defparam i1145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1144_3_lut (.I0(ram_s_63_0), .I1(register_vector[8]), .I2(n194), 
            .I3(GND_net), .O(n1392));   // src/ram.vhd(56[12:17])
    defparam i1144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1143_3_lut (.I0(ram_s_62_7), .I1(sx[7]), .I2(n195), .I3(GND_net), 
            .O(n1391));   // src/ram.vhd(56[12:17])
    defparam i1143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1142_3_lut (.I0(ram_s_62_6), .I1(sx[6]), .I2(n195), .I3(GND_net), 
            .O(n1390));   // src/ram.vhd(56[12:17])
    defparam i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1141_3_lut (.I0(ram_s_62_5), .I1(sx[5]), .I2(n195), .I3(GND_net), 
            .O(n1389));   // src/ram.vhd(56[12:17])
    defparam i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1140_3_lut (.I0(ram_s_62_4), .I1(sx[4]), .I2(n195), .I3(GND_net), 
            .O(n1388));   // src/ram.vhd(56[12:17])
    defparam i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1139_3_lut (.I0(ram_s_62_3), .I1(register_vector[11]), .I2(n195), 
            .I3(GND_net), .O(n1387));   // src/ram.vhd(56[12:17])
    defparam i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1138_3_lut (.I0(ram_s_62_2), .I1(register_vector[10]), .I2(n195), 
            .I3(GND_net), .O(n1386));   // src/ram.vhd(56[12:17])
    defparam i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1137_3_lut (.I0(ram_s_62_1), .I1(register_vector[9]), .I2(n195), 
            .I3(GND_net), .O(n1385));   // src/ram.vhd(56[12:17])
    defparam i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1136_3_lut (.I0(ram_s_62_0), .I1(register_vector[8]), .I2(n195), 
            .I3(GND_net), .O(n1384));   // src/ram.vhd(56[12:17])
    defparam i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1111_3_lut (.I0(ram_s_58_7), .I1(sx[7]), .I2(n199), .I3(GND_net), 
            .O(n1359));   // src/ram.vhd(56[12:17])
    defparam i1111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1110_3_lut (.I0(ram_s_58_6), .I1(sx[6]), .I2(n199), .I3(GND_net), 
            .O(n1358));   // src/ram.vhd(56[12:17])
    defparam i1110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1109_3_lut (.I0(ram_s_58_5), .I1(sx[5]), .I2(n199), .I3(GND_net), 
            .O(n1357));   // src/ram.vhd(56[12:17])
    defparam i1109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1108_3_lut (.I0(ram_s_58_4), .I1(sx[4]), .I2(n199), .I3(GND_net), 
            .O(n1356));   // src/ram.vhd(56[12:17])
    defparam i1108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1107_3_lut (.I0(ram_s_58_3), .I1(register_vector[11]), .I2(n199), 
            .I3(GND_net), .O(n1355));   // src/ram.vhd(56[12:17])
    defparam i1107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1106_3_lut (.I0(ram_s_58_2), .I1(register_vector[10]), .I2(n199), 
            .I3(GND_net), .O(n1354));   // src/ram.vhd(56[12:17])
    defparam i1106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1105_3_lut (.I0(ram_s_58_1), .I1(register_vector[9]), .I2(n199), 
            .I3(GND_net), .O(n1353));   // src/ram.vhd(56[12:17])
    defparam i1105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1104_3_lut (.I0(ram_s_58_0), .I1(register_vector[8]), .I2(n199), 
            .I3(GND_net), .O(n1352));   // src/ram.vhd(56[12:17])
    defparam i1104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1103_3_lut (.I0(ram_s_57_7), .I1(sx[7]), .I2(n200), .I3(GND_net), 
            .O(n1351));   // src/ram.vhd(56[12:17])
    defparam i1103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1102_3_lut (.I0(ram_s_57_6), .I1(sx[6]), .I2(n200), .I3(GND_net), 
            .O(n1350));   // src/ram.vhd(56[12:17])
    defparam i1102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1101_3_lut (.I0(ram_s_57_5), .I1(sx[5]), .I2(n200), .I3(GND_net), 
            .O(n1349));   // src/ram.vhd(56[12:17])
    defparam i1101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1100_3_lut (.I0(ram_s_57_4), .I1(sx[4]), .I2(n200), .I3(GND_net), 
            .O(n1348));   // src/ram.vhd(56[12:17])
    defparam i1100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1099_3_lut (.I0(ram_s_57_3), .I1(register_vector[11]), .I2(n200), 
            .I3(GND_net), .O(n1347));   // src/ram.vhd(56[12:17])
    defparam i1099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1098_3_lut (.I0(ram_s_57_2), .I1(register_vector[10]), .I2(n200), 
            .I3(GND_net), .O(n1346));   // src/ram.vhd(56[12:17])
    defparam i1098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1097_3_lut (.I0(ram_s_57_1), .I1(register_vector[9]), .I2(n200), 
            .I3(GND_net), .O(n1345));   // src/ram.vhd(56[12:17])
    defparam i1097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1096_3_lut (.I0(ram_s_57_0), .I1(register_vector[8]), .I2(n200), 
            .I3(GND_net), .O(n1344));   // src/ram.vhd(56[12:17])
    defparam i1096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1023_3_lut (.I0(ram_s_47_7), .I1(sx[7]), .I2(n210), .I3(GND_net), 
            .O(n1271));   // src/ram.vhd(56[12:17])
    defparam i1023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1022_3_lut (.I0(ram_s_47_6), .I1(sx[6]), .I2(n210), .I3(GND_net), 
            .O(n1270));   // src/ram.vhd(56[12:17])
    defparam i1022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1021_3_lut (.I0(ram_s_47_5), .I1(sx[5]), .I2(n210), .I3(GND_net), 
            .O(n1269));   // src/ram.vhd(56[12:17])
    defparam i1021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1020_3_lut (.I0(ram_s_47_4), .I1(sx[4]), .I2(n210), .I3(GND_net), 
            .O(n1268));   // src/ram.vhd(56[12:17])
    defparam i1020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1019_3_lut (.I0(ram_s_47_3), .I1(register_vector[11]), .I2(n210), 
            .I3(GND_net), .O(n1267));   // src/ram.vhd(56[12:17])
    defparam i1019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1018_3_lut (.I0(ram_s_47_2), .I1(register_vector[10]), .I2(n210), 
            .I3(GND_net), .O(n1266));   // src/ram.vhd(56[12:17])
    defparam i1018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1017_3_lut (.I0(ram_s_47_1), .I1(register_vector[9]), .I2(n210), 
            .I3(GND_net), .O(n1265));   // src/ram.vhd(56[12:17])
    defparam i1017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1016_3_lut (.I0(ram_s_47_0), .I1(register_vector[8]), .I2(n210), 
            .I3(GND_net), .O(n1264));   // src/ram.vhd(56[12:17])
    defparam i1016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1007_3_lut (.I0(ram_s_45_7), .I1(sx[7]), .I2(n212), .I3(GND_net), 
            .O(n1255));   // src/ram.vhd(56[12:17])
    defparam i1007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1006_3_lut (.I0(ram_s_45_6), .I1(sx[6]), .I2(n212), .I3(GND_net), 
            .O(n1254));   // src/ram.vhd(56[12:17])
    defparam i1006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1005_3_lut (.I0(ram_s_45_5), .I1(sx[5]), .I2(n212), .I3(GND_net), 
            .O(n1253));   // src/ram.vhd(56[12:17])
    defparam i1005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1004_3_lut (.I0(ram_s_45_4), .I1(sx[4]), .I2(n212), .I3(GND_net), 
            .O(n1252));   // src/ram.vhd(56[12:17])
    defparam i1004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1003_3_lut (.I0(ram_s_45_3), .I1(register_vector[11]), .I2(n212), 
            .I3(GND_net), .O(n1251));   // src/ram.vhd(56[12:17])
    defparam i1003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1002_3_lut (.I0(ram_s_45_2), .I1(register_vector[10]), .I2(n212), 
            .I3(GND_net), .O(n1250));   // src/ram.vhd(56[12:17])
    defparam i1002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1001_3_lut (.I0(ram_s_45_1), .I1(register_vector[9]), .I2(n212), 
            .I3(GND_net), .O(n1249));   // src/ram.vhd(56[12:17])
    defparam i1001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1000_3_lut (.I0(ram_s_45_0), .I1(register_vector[8]), .I2(n212), 
            .I3(GND_net), .O(n1248));   // src/ram.vhd(56[12:17])
    defparam i1000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i999_3_lut (.I0(ram_s_44_7), .I1(sx[7]), .I2(n213), .I3(GND_net), 
            .O(n1247));   // src/ram.vhd(56[12:17])
    defparam i999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i998_3_lut (.I0(ram_s_44_6), .I1(sx[6]), .I2(n213), .I3(GND_net), 
            .O(n1246));   // src/ram.vhd(56[12:17])
    defparam i998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i997_3_lut (.I0(ram_s_44_5), .I1(sx[5]), .I2(n213), .I3(GND_net), 
            .O(n1245));   // src/ram.vhd(56[12:17])
    defparam i997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i996_3_lut (.I0(ram_s_44_4), .I1(sx[4]), .I2(n213), .I3(GND_net), 
            .O(n1244));   // src/ram.vhd(56[12:17])
    defparam i996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i995_3_lut (.I0(ram_s_44_3), .I1(register_vector[11]), .I2(n213), 
            .I3(GND_net), .O(n1243));   // src/ram.vhd(56[12:17])
    defparam i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i994_3_lut (.I0(ram_s_44_2), .I1(register_vector[10]), .I2(n213), 
            .I3(GND_net), .O(n1242));   // src/ram.vhd(56[12:17])
    defparam i994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i993_3_lut (.I0(ram_s_44_1), .I1(register_vector[9]), .I2(n213), 
            .I3(GND_net), .O(n1241));   // src/ram.vhd(56[12:17])
    defparam i993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i992_3_lut (.I0(ram_s_44_0), .I1(register_vector[8]), .I2(n213), 
            .I3(GND_net), .O(n1240));   // src/ram.vhd(56[12:17])
    defparam i992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i991_3_lut (.I0(ram_s_43_7), .I1(sx[7]), .I2(n214), .I3(GND_net), 
            .O(n1239));   // src/ram.vhd(56[12:17])
    defparam i991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i990_3_lut (.I0(ram_s_43_6), .I1(sx[6]), .I2(n214), .I3(GND_net), 
            .O(n1238));   // src/ram.vhd(56[12:17])
    defparam i990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i989_3_lut (.I0(ram_s_43_5), .I1(sx[5]), .I2(n214), .I3(GND_net), 
            .O(n1237));   // src/ram.vhd(56[12:17])
    defparam i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i988_3_lut (.I0(ram_s_43_4), .I1(sx[4]), .I2(n214), .I3(GND_net), 
            .O(n1236));   // src/ram.vhd(56[12:17])
    defparam i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i987_3_lut (.I0(ram_s_43_3), .I1(register_vector[11]), .I2(n214), 
            .I3(GND_net), .O(n1235));   // src/ram.vhd(56[12:17])
    defparam i987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i986_3_lut (.I0(ram_s_43_2), .I1(register_vector[10]), .I2(n214), 
            .I3(GND_net), .O(n1234));   // src/ram.vhd(56[12:17])
    defparam i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i985_3_lut (.I0(ram_s_43_1), .I1(register_vector[9]), .I2(n214), 
            .I3(GND_net), .O(n1233));   // src/ram.vhd(56[12:17])
    defparam i985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i984_3_lut (.I0(ram_s_43_0), .I1(register_vector[8]), .I2(n214), 
            .I3(GND_net), .O(n1232));   // src/ram.vhd(56[12:17])
    defparam i984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i967_3_lut (.I0(ram_s_40_7), .I1(sx[7]), .I2(n217), .I3(GND_net), 
            .O(n1215));   // src/ram.vhd(56[12:17])
    defparam i967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i966_3_lut (.I0(ram_s_40_6), .I1(sx[6]), .I2(n217), .I3(GND_net), 
            .O(n1214));   // src/ram.vhd(56[12:17])
    defparam i966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i965_3_lut (.I0(ram_s_40_5), .I1(sx[5]), .I2(n217), .I3(GND_net), 
            .O(n1213));   // src/ram.vhd(56[12:17])
    defparam i965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i964_3_lut (.I0(ram_s_40_4), .I1(sx[4]), .I2(n217), .I3(GND_net), 
            .O(n1212));   // src/ram.vhd(56[12:17])
    defparam i964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i963_3_lut (.I0(ram_s_40_3), .I1(register_vector[11]), .I2(n217), 
            .I3(GND_net), .O(n1211));   // src/ram.vhd(56[12:17])
    defparam i963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i962_3_lut (.I0(ram_s_40_2), .I1(register_vector[10]), .I2(n217), 
            .I3(GND_net), .O(n1210));   // src/ram.vhd(56[12:17])
    defparam i962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i961_3_lut (.I0(ram_s_40_1), .I1(register_vector[9]), .I2(n217), 
            .I3(GND_net), .O(n1209));   // src/ram.vhd(56[12:17])
    defparam i961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i960_3_lut (.I0(ram_s_40_0), .I1(register_vector[8]), .I2(n217), 
            .I3(GND_net), .O(n1208));   // src/ram.vhd(56[12:17])
    defparam i960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i959_3_lut (.I0(ram_s_39_7), .I1(sx[7]), .I2(n218), .I3(GND_net), 
            .O(n1207));   // src/ram.vhd(56[12:17])
    defparam i959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i958_3_lut (.I0(ram_s_39_6), .I1(sx[6]), .I2(n218), .I3(GND_net), 
            .O(n1206));   // src/ram.vhd(56[12:17])
    defparam i958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i957_3_lut (.I0(ram_s_39_5), .I1(sx[5]), .I2(n218), .I3(GND_net), 
            .O(n1205));   // src/ram.vhd(56[12:17])
    defparam i957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i956_3_lut (.I0(ram_s_39_4), .I1(sx[4]), .I2(n218), .I3(GND_net), 
            .O(n1204));   // src/ram.vhd(56[12:17])
    defparam i956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i955_3_lut (.I0(ram_s_39_3), .I1(register_vector[11]), .I2(n218), 
            .I3(GND_net), .O(n1203));   // src/ram.vhd(56[12:17])
    defparam i955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i954_3_lut (.I0(ram_s_39_2), .I1(register_vector[10]), .I2(n218), 
            .I3(GND_net), .O(n1202));   // src/ram.vhd(56[12:17])
    defparam i954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i953_3_lut (.I0(ram_s_39_1), .I1(register_vector[9]), .I2(n218), 
            .I3(GND_net), .O(n1201));   // src/ram.vhd(56[12:17])
    defparam i953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i952_3_lut (.I0(ram_s_39_0), .I1(register_vector[8]), .I2(n218), 
            .I3(GND_net), .O(n1200));   // src/ram.vhd(56[12:17])
    defparam i952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i951_3_lut (.I0(ram_s_38_7), .I1(sx[7]), .I2(n219), .I3(GND_net), 
            .O(n1199));   // src/ram.vhd(56[12:17])
    defparam i951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i950_3_lut (.I0(ram_s_38_6), .I1(sx[6]), .I2(n219), .I3(GND_net), 
            .O(n1198));   // src/ram.vhd(56[12:17])
    defparam i950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i949_3_lut (.I0(ram_s_38_5), .I1(sx[5]), .I2(n219), .I3(GND_net), 
            .O(n1197));   // src/ram.vhd(56[12:17])
    defparam i949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i948_3_lut (.I0(ram_s_38_4), .I1(sx[4]), .I2(n219), .I3(GND_net), 
            .O(n1196));   // src/ram.vhd(56[12:17])
    defparam i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i947_3_lut (.I0(ram_s_38_3), .I1(register_vector[11]), .I2(n219), 
            .I3(GND_net), .O(n1195));   // src/ram.vhd(56[12:17])
    defparam i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i946_3_lut (.I0(ram_s_38_2), .I1(register_vector[10]), .I2(n219), 
            .I3(GND_net), .O(n1194));   // src/ram.vhd(56[12:17])
    defparam i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i945_3_lut (.I0(ram_s_38_1), .I1(register_vector[9]), .I2(n219), 
            .I3(GND_net), .O(n1193));   // src/ram.vhd(56[12:17])
    defparam i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i944_3_lut (.I0(ram_s_38_0), .I1(register_vector[8]), .I2(n219), 
            .I3(GND_net), .O(n1192));   // src/ram.vhd(56[12:17])
    defparam i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i943_3_lut (.I0(ram_s_37_7), .I1(sx[7]), .I2(n220), .I3(GND_net), 
            .O(n1191));   // src/ram.vhd(56[12:17])
    defparam i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i942_3_lut (.I0(ram_s_37_6), .I1(sx[6]), .I2(n220), .I3(GND_net), 
            .O(n1190));   // src/ram.vhd(56[12:17])
    defparam i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i941_3_lut (.I0(ram_s_37_5), .I1(sx[5]), .I2(n220), .I3(GND_net), 
            .O(n1189));   // src/ram.vhd(56[12:17])
    defparam i941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i940_3_lut (.I0(ram_s_37_4), .I1(sx[4]), .I2(n220), .I3(GND_net), 
            .O(n1188));   // src/ram.vhd(56[12:17])
    defparam i940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i939_3_lut (.I0(ram_s_37_3), .I1(register_vector[11]), .I2(n220), 
            .I3(GND_net), .O(n1187));   // src/ram.vhd(56[12:17])
    defparam i939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i938_3_lut (.I0(ram_s_37_2), .I1(register_vector[10]), .I2(n220), 
            .I3(GND_net), .O(n1186));   // src/ram.vhd(56[12:17])
    defparam i938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i937_3_lut (.I0(ram_s_37_1), .I1(register_vector[9]), .I2(n220), 
            .I3(GND_net), .O(n1185));   // src/ram.vhd(56[12:17])
    defparam i937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i936_3_lut (.I0(ram_s_37_0), .I1(register_vector[8]), .I2(n220), 
            .I3(GND_net), .O(n1184));   // src/ram.vhd(56[12:17])
    defparam i936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i935_3_lut (.I0(ram_s_36_7), .I1(sx[7]), .I2(n221), .I3(GND_net), 
            .O(n1183));   // src/ram.vhd(56[12:17])
    defparam i935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i934_3_lut (.I0(ram_s_36_6), .I1(sx[6]), .I2(n221), .I3(GND_net), 
            .O(n1182));   // src/ram.vhd(56[12:17])
    defparam i934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i933_3_lut (.I0(ram_s_36_5), .I1(sx[5]), .I2(n221), .I3(GND_net), 
            .O(n1181));   // src/ram.vhd(56[12:17])
    defparam i933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i932_3_lut (.I0(ram_s_36_4), .I1(sx[4]), .I2(n221), .I3(GND_net), 
            .O(n1180));   // src/ram.vhd(56[12:17])
    defparam i932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i931_3_lut (.I0(ram_s_36_3), .I1(register_vector[11]), .I2(n221), 
            .I3(GND_net), .O(n1179));   // src/ram.vhd(56[12:17])
    defparam i931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i930_3_lut (.I0(ram_s_36_2), .I1(register_vector[10]), .I2(n221), 
            .I3(GND_net), .O(n1178));   // src/ram.vhd(56[12:17])
    defparam i930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i929_3_lut (.I0(ram_s_36_1), .I1(register_vector[9]), .I2(n221), 
            .I3(GND_net), .O(n1177));   // src/ram.vhd(56[12:17])
    defparam i929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i928_3_lut (.I0(ram_s_36_0), .I1(register_vector[8]), .I2(n221), 
            .I3(GND_net), .O(n1176));   // src/ram.vhd(56[12:17])
    defparam i928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i927_3_lut (.I0(ram_s_35_7), .I1(sx[7]), .I2(n222), .I3(GND_net), 
            .O(n1175));   // src/ram.vhd(56[12:17])
    defparam i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i926_3_lut (.I0(ram_s_35_6), .I1(sx[6]), .I2(n222), .I3(GND_net), 
            .O(n1174));   // src/ram.vhd(56[12:17])
    defparam i926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i925_3_lut (.I0(ram_s_35_5), .I1(sx[5]), .I2(n222), .I3(GND_net), 
            .O(n1173));   // src/ram.vhd(56[12:17])
    defparam i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i924_3_lut (.I0(ram_s_35_4), .I1(sx[4]), .I2(n222), .I3(GND_net), 
            .O(n1172));   // src/ram.vhd(56[12:17])
    defparam i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i923_3_lut (.I0(ram_s_35_3), .I1(register_vector[11]), .I2(n222), 
            .I3(GND_net), .O(n1171));   // src/ram.vhd(56[12:17])
    defparam i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i922_3_lut (.I0(ram_s_35_2), .I1(register_vector[10]), .I2(n222), 
            .I3(GND_net), .O(n1170));   // src/ram.vhd(56[12:17])
    defparam i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i921_3_lut (.I0(ram_s_35_1), .I1(register_vector[9]), .I2(n222), 
            .I3(GND_net), .O(n1169));   // src/ram.vhd(56[12:17])
    defparam i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i920_3_lut (.I0(ram_s_35_0), .I1(register_vector[8]), .I2(n222), 
            .I3(GND_net), .O(n1168));   // src/ram.vhd(56[12:17])
    defparam i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i919_3_lut (.I0(ram_s_34_7), .I1(sx[7]), .I2(n223), .I3(GND_net), 
            .O(n1167));   // src/ram.vhd(56[12:17])
    defparam i919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i918_3_lut (.I0(ram_s_34_6), .I1(sx[6]), .I2(n223), .I3(GND_net), 
            .O(n1166));   // src/ram.vhd(56[12:17])
    defparam i918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i917_3_lut (.I0(ram_s_34_5), .I1(sx[5]), .I2(n223), .I3(GND_net), 
            .O(n1165));   // src/ram.vhd(56[12:17])
    defparam i917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i916_3_lut (.I0(ram_s_34_4), .I1(sx[4]), .I2(n223), .I3(GND_net), 
            .O(n1164));   // src/ram.vhd(56[12:17])
    defparam i916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i915_3_lut (.I0(ram_s_34_3), .I1(register_vector[11]), .I2(n223), 
            .I3(GND_net), .O(n1163));   // src/ram.vhd(56[12:17])
    defparam i915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i914_3_lut (.I0(ram_s_34_2), .I1(register_vector[10]), .I2(n223), 
            .I3(GND_net), .O(n1162));   // src/ram.vhd(56[12:17])
    defparam i914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i913_3_lut (.I0(ram_s_34_1), .I1(register_vector[9]), .I2(n223), 
            .I3(GND_net), .O(n1161));   // src/ram.vhd(56[12:17])
    defparam i913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i912_3_lut (.I0(ram_s_34_0), .I1(register_vector[8]), .I2(n223), 
            .I3(GND_net), .O(n1160));   // src/ram.vhd(56[12:17])
    defparam i912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i911_3_lut (.I0(ram_s_33_7), .I1(sx[7]), .I2(n224), .I3(GND_net), 
            .O(n1159));   // src/ram.vhd(56[12:17])
    defparam i911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i910_3_lut (.I0(ram_s_33_6), .I1(sx[6]), .I2(n224), .I3(GND_net), 
            .O(n1158));   // src/ram.vhd(56[12:17])
    defparam i910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i909_3_lut (.I0(ram_s_33_5), .I1(sx[5]), .I2(n224), .I3(GND_net), 
            .O(n1157));   // src/ram.vhd(56[12:17])
    defparam i909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i908_3_lut (.I0(ram_s_33_4), .I1(sx[4]), .I2(n224), .I3(GND_net), 
            .O(n1156));   // src/ram.vhd(56[12:17])
    defparam i908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i907_3_lut (.I0(ram_s_33_3), .I1(register_vector[11]), .I2(n224), 
            .I3(GND_net), .O(n1155));   // src/ram.vhd(56[12:17])
    defparam i907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i906_3_lut (.I0(ram_s_33_2), .I1(register_vector[10]), .I2(n224), 
            .I3(GND_net), .O(n1154));   // src/ram.vhd(56[12:17])
    defparam i906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i905_3_lut (.I0(ram_s_33_1), .I1(register_vector[9]), .I2(n224), 
            .I3(GND_net), .O(n1153));   // src/ram.vhd(56[12:17])
    defparam i905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i904_3_lut (.I0(ram_s_33_0), .I1(register_vector[8]), .I2(n224), 
            .I3(GND_net), .O(n1152));   // src/ram.vhd(56[12:17])
    defparam i904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i903_3_lut (.I0(ram_s_32_7), .I1(sx[7]), .I2(n225), .I3(GND_net), 
            .O(n1151));   // src/ram.vhd(56[12:17])
    defparam i903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i902_3_lut (.I0(ram_s_32_6), .I1(sx[6]), .I2(n225), .I3(GND_net), 
            .O(n1150));   // src/ram.vhd(56[12:17])
    defparam i902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i901_3_lut (.I0(ram_s_32_5), .I1(sx[5]), .I2(n225), .I3(GND_net), 
            .O(n1149));   // src/ram.vhd(56[12:17])
    defparam i901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i900_3_lut (.I0(ram_s_32_4), .I1(sx[4]), .I2(n225), .I3(GND_net), 
            .O(n1148));   // src/ram.vhd(56[12:17])
    defparam i900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i899_3_lut (.I0(ram_s_32_3), .I1(register_vector[11]), .I2(n225), 
            .I3(GND_net), .O(n1147));   // src/ram.vhd(56[12:17])
    defparam i899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i898_3_lut (.I0(ram_s_32_2), .I1(register_vector[10]), .I2(n225), 
            .I3(GND_net), .O(n1146));   // src/ram.vhd(56[12:17])
    defparam i898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i897_3_lut (.I0(ram_s_32_1), .I1(register_vector[9]), .I2(n225), 
            .I3(GND_net), .O(n1145));   // src/ram.vhd(56[12:17])
    defparam i897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i896_3_lut (.I0(ram_s_32_0), .I1(register_vector[8]), .I2(n225), 
            .I3(GND_net), .O(n1144));   // src/ram.vhd(56[12:17])
    defparam i896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i803_3_lut (.I0(ram_s_14_5), .I1(sx[5]), .I2(n243), .I3(GND_net), 
            .O(n1051));   // src/ram.vhd(56[12:17])
    defparam i803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i799_3_lut (.I0(ram_s_0_0), .I1(register_vector[8]), .I2(n257), 
            .I3(GND_net), .O(n1047));   // src/ram.vhd(56[12:17])
    defparam i799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i798_3_lut (.I0(ram_s_0_1), .I1(register_vector[9]), .I2(n257), 
            .I3(GND_net), .O(n1046));   // src/ram.vhd(56[12:17])
    defparam i798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i797_3_lut (.I0(ram_s_0_2), .I1(register_vector[10]), .I2(n257), 
            .I3(GND_net), .O(n1045));   // src/ram.vhd(56[12:17])
    defparam i797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i796_3_lut (.I0(ram_s_12_3), .I1(register_vector[11]), .I2(n245), 
            .I3(GND_net), .O(n1044));   // src/ram.vhd(56[12:17])
    defparam i796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i795_3_lut (.I0(ram_s_11_6), .I1(sx[6]), .I2(n246), .I3(GND_net), 
            .O(n1043));   // src/ram.vhd(56[12:17])
    defparam i795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i794_3_lut (.I0(ram_s_11_1), .I1(register_vector[9]), .I2(n246), 
            .I3(GND_net), .O(n1042));   // src/ram.vhd(56[12:17])
    defparam i794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i793_3_lut (.I0(ram_s_12_6), .I1(sx[6]), .I2(n245), .I3(GND_net), 
            .O(n1041));   // src/ram.vhd(56[12:17])
    defparam i793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i792_3_lut (.I0(ram_s_12_1), .I1(register_vector[9]), .I2(n245), 
            .I3(GND_net), .O(n1040));   // src/ram.vhd(56[12:17])
    defparam i792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i790_3_lut (.I0(ram_s_11_4), .I1(sx[4]), .I2(n246), .I3(GND_net), 
            .O(n1038));   // src/ram.vhd(56[12:17])
    defparam i790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i789_3_lut (.I0(ram_s_12_4), .I1(sx[4]), .I2(n245), .I3(GND_net), 
            .O(n1037));   // src/ram.vhd(56[12:17])
    defparam i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i788_3_lut (.I0(ram_s_11_7), .I1(sx[7]), .I2(n246), .I3(GND_net), 
            .O(n1036));   // src/ram.vhd(56[12:17])
    defparam i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i787_3_lut (.I0(ram_s_11_2), .I1(register_vector[10]), .I2(n246), 
            .I3(GND_net), .O(n1035));   // src/ram.vhd(56[12:17])
    defparam i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i786_3_lut (.I0(ram_s_12_7), .I1(sx[7]), .I2(n245), .I3(GND_net), 
            .O(n1034));   // src/ram.vhd(56[12:17])
    defparam i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i785_3_lut (.I0(ram_s_12_2), .I1(register_vector[10]), .I2(n245), 
            .I3(GND_net), .O(n1033));   // src/ram.vhd(56[12:17])
    defparam i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i784_3_lut (.I0(ram_s_11_5), .I1(sx[5]), .I2(n246), .I3(GND_net), 
            .O(n1032));   // src/ram.vhd(56[12:17])
    defparam i784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i783_3_lut (.I0(ram_s_12_5), .I1(sx[5]), .I2(n245), .I3(GND_net), 
            .O(n1031));   // src/ram.vhd(56[12:17])
    defparam i783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i782_3_lut (.I0(ram_s_12_0), .I1(register_vector[8]), .I2(n245), 
            .I3(GND_net), .O(n1030));   // src/ram.vhd(56[12:17])
    defparam i782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i781_3_lut (.I0(ram_s_11_3), .I1(register_vector[11]), .I2(n246), 
            .I3(GND_net), .O(n1029));   // src/ram.vhd(56[12:17])
    defparam i781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i769_3_lut (.I0(ram_s_0_3), .I1(register_vector[11]), .I2(n257), 
            .I3(GND_net), .O(n1017));   // src/ram.vhd(56[12:17])
    defparam i769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i768_3_lut (.I0(ram_s_0_4), .I1(sx[4]), .I2(n257), .I3(GND_net), 
            .O(n1016));   // src/ram.vhd(56[12:17])
    defparam i768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i767_3_lut (.I0(ram_s_0_5), .I1(sx[5]), .I2(n257), .I3(GND_net), 
            .O(n1015));   // src/ram.vhd(56[12:17])
    defparam i767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i766_3_lut (.I0(ram_s_0_6), .I1(sx[6]), .I2(n257), .I3(GND_net), 
            .O(n1014));   // src/ram.vhd(56[12:17])
    defparam i766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i765_3_lut (.I0(ram_s_0_7), .I1(sx[7]), .I2(n257), .I3(GND_net), 
            .O(n1013));   // src/ram.vhd(56[12:17])
    defparam i765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i764_3_lut (.I0(ram_s_1_0), .I1(register_vector[8]), .I2(n256), 
            .I3(GND_net), .O(n1012));   // src/ram.vhd(56[12:17])
    defparam i764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i763_3_lut (.I0(ram_s_1_1), .I1(register_vector[9]), .I2(n256), 
            .I3(GND_net), .O(n1011));   // src/ram.vhd(56[12:17])
    defparam i763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i762_3_lut (.I0(ram_s_1_2), .I1(register_vector[10]), .I2(n256), 
            .I3(GND_net), .O(n1010));   // src/ram.vhd(56[12:17])
    defparam i762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i761_3_lut (.I0(ram_s_1_3), .I1(register_vector[11]), .I2(n256), 
            .I3(GND_net), .O(n1009));   // src/ram.vhd(56[12:17])
    defparam i761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i760_3_lut (.I0(ram_s_1_4), .I1(sx[4]), .I2(n256), .I3(GND_net), 
            .O(n1008));   // src/ram.vhd(56[12:17])
    defparam i760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i759_3_lut (.I0(ram_s_1_5), .I1(sx[5]), .I2(n256), .I3(GND_net), 
            .O(n1007));   // src/ram.vhd(56[12:17])
    defparam i759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i758_3_lut (.I0(ram_s_4_4), .I1(sx[4]), .I2(n253), .I3(GND_net), 
            .O(n1006));   // src/ram.vhd(56[12:17])
    defparam i758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i757_3_lut (.I0(ram_s_4_7), .I1(sx[7]), .I2(n253), .I3(GND_net), 
            .O(n1005));   // src/ram.vhd(56[12:17])
    defparam i757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i756_3_lut (.I0(ram_s_4_5), .I1(sx[5]), .I2(n253), .I3(GND_net), 
            .O(n1004));   // src/ram.vhd(56[12:17])
    defparam i756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i755_3_lut (.I0(ram_s_5_0), .I1(register_vector[8]), .I2(n252), 
            .I3(GND_net), .O(n1003));   // src/ram.vhd(56[12:17])
    defparam i755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i754_3_lut (.I0(ram_s_4_6), .I1(sx[6]), .I2(n253), .I3(GND_net), 
            .O(n1002));   // src/ram.vhd(56[12:17])
    defparam i754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i753_3_lut (.I0(ram_s_5_1), .I1(register_vector[9]), .I2(n252), 
            .I3(GND_net), .O(n1001));   // src/ram.vhd(56[12:17])
    defparam i753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i750_3_lut (.I0(ram_s_8_5), .I1(sx[5]), .I2(n249), .I3(GND_net), 
            .O(n998));   // src/ram.vhd(56[12:17])
    defparam i750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i749_3_lut (.I0(ram_s_8_2), .I1(register_vector[10]), .I2(n249), 
            .I3(GND_net), .O(n997));   // src/ram.vhd(56[12:17])
    defparam i749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i748_3_lut (.I0(ram_s_7_7), .I1(sx[7]), .I2(n250), .I3(GND_net), 
            .O(n996));   // src/ram.vhd(56[12:17])
    defparam i748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i747_3_lut (.I0(ram_s_7_4), .I1(sx[4]), .I2(n250), .I3(GND_net), 
            .O(n995));   // src/ram.vhd(56[12:17])
    defparam i747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i746_3_lut (.I0(ram_s_7_1), .I1(register_vector[9]), .I2(n250), 
            .I3(GND_net), .O(n994));   // src/ram.vhd(56[12:17])
    defparam i746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i745_3_lut (.I0(ram_s_6_6), .I1(sx[6]), .I2(n251), .I3(GND_net), 
            .O(n993));   // src/ram.vhd(56[12:17])
    defparam i745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i744_3_lut (.I0(ram_s_6_3), .I1(register_vector[11]), .I2(n251), 
            .I3(GND_net), .O(n992));   // src/ram.vhd(56[12:17])
    defparam i744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i741_3_lut (.I0(ram_s_8_6), .I1(sx[6]), .I2(n249), .I3(GND_net), 
            .O(n989));   // src/ram.vhd(56[12:17])
    defparam i741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i740_3_lut (.I0(ram_s_8_3), .I1(register_vector[11]), .I2(n249), 
            .I3(GND_net), .O(n988));   // src/ram.vhd(56[12:17])
    defparam i740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i739_3_lut (.I0(ram_s_8_0), .I1(register_vector[8]), .I2(n249), 
            .I3(GND_net), .O(n987));   // src/ram.vhd(56[12:17])
    defparam i739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i738_3_lut (.I0(ram_s_7_5), .I1(sx[5]), .I2(n250), .I3(GND_net), 
            .O(n986));   // src/ram.vhd(56[12:17])
    defparam i738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i737_3_lut (.I0(ram_s_7_2), .I1(register_vector[10]), .I2(n250), 
            .I3(GND_net), .O(n985));   // src/ram.vhd(56[12:17])
    defparam i737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i736_3_lut (.I0(ram_s_6_7), .I1(sx[7]), .I2(n251), .I3(GND_net), 
            .O(n984));   // src/ram.vhd(56[12:17])
    defparam i736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i735_3_lut (.I0(ram_s_6_4), .I1(sx[4]), .I2(n251), .I3(GND_net), 
            .O(n983));   // src/ram.vhd(56[12:17])
    defparam i735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i732_3_lut (.I0(ram_s_8_7), .I1(sx[7]), .I2(n249), .I3(GND_net), 
            .O(n980));   // src/ram.vhd(56[12:17])
    defparam i732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i731_3_lut (.I0(ram_s_8_4), .I1(sx[4]), .I2(n249), .I3(GND_net), 
            .O(n979));   // src/ram.vhd(56[12:17])
    defparam i731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i730_3_lut (.I0(ram_s_8_1), .I1(register_vector[9]), .I2(n249), 
            .I3(GND_net), .O(n978));   // src/ram.vhd(56[12:17])
    defparam i730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i729_3_lut (.I0(ram_s_7_6), .I1(sx[6]), .I2(n250), .I3(GND_net), 
            .O(n977));   // src/ram.vhd(56[12:17])
    defparam i729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i728_3_lut (.I0(ram_s_7_3), .I1(register_vector[11]), .I2(n250), 
            .I3(GND_net), .O(n976));   // src/ram.vhd(56[12:17])
    defparam i728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i727_3_lut (.I0(ram_s_7_0), .I1(register_vector[8]), .I2(n250), 
            .I3(GND_net), .O(n975));   // src/ram.vhd(56[12:17])
    defparam i727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i726_3_lut (.I0(ram_s_6_5), .I1(sx[5]), .I2(n251), .I3(GND_net), 
            .O(n974));   // src/ram.vhd(56[12:17])
    defparam i726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i725_3_lut (.I0(ram_s_1_6), .I1(sx[6]), .I2(n256), .I3(GND_net), 
            .O(n973));   // src/ram.vhd(56[12:17])
    defparam i725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i724_3_lut (.I0(ram_s_1_7), .I1(sx[7]), .I2(n256), .I3(GND_net), 
            .O(n972));   // src/ram.vhd(56[12:17])
    defparam i724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i723_3_lut (.I0(ram_s_2_0), .I1(register_vector[8]), .I2(n255), 
            .I3(GND_net), .O(n971));   // src/ram.vhd(56[12:17])
    defparam i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i722_3_lut (.I0(ram_s_2_1), .I1(register_vector[9]), .I2(n255), 
            .I3(GND_net), .O(n970));   // src/ram.vhd(56[12:17])
    defparam i722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i721_3_lut (.I0(ram_s_2_2), .I1(register_vector[10]), .I2(n255), 
            .I3(GND_net), .O(n969));   // src/ram.vhd(56[12:17])
    defparam i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i720_3_lut (.I0(ram_s_2_3), .I1(register_vector[11]), .I2(n255), 
            .I3(GND_net), .O(n968));   // src/ram.vhd(56[12:17])
    defparam i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i719_3_lut (.I0(ram_s_2_4), .I1(sx[4]), .I2(n255), .I3(GND_net), 
            .O(n967));   // src/ram.vhd(56[12:17])
    defparam i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i718_3_lut (.I0(ram_s_2_5), .I1(sx[5]), .I2(n255), .I3(GND_net), 
            .O(n966));   // src/ram.vhd(56[12:17])
    defparam i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i717_3_lut (.I0(ram_s_2_6), .I1(sx[6]), .I2(n255), .I3(GND_net), 
            .O(n965));   // src/ram.vhd(56[12:17])
    defparam i717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i716_3_lut (.I0(ram_s_2_7), .I1(sx[7]), .I2(n255), .I3(GND_net), 
            .O(n964));   // src/ram.vhd(56[12:17])
    defparam i716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i715_3_lut (.I0(ram_s_3_0), .I1(register_vector[8]), .I2(n254), 
            .I3(GND_net), .O(n963));   // src/ram.vhd(56[12:17])
    defparam i715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i714_3_lut (.I0(ram_s_3_1), .I1(register_vector[9]), .I2(n254), 
            .I3(GND_net), .O(n962));   // src/ram.vhd(56[12:17])
    defparam i714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i713_3_lut (.I0(ram_s_3_2), .I1(register_vector[10]), .I2(n254), 
            .I3(GND_net), .O(n961));   // src/ram.vhd(56[12:17])
    defparam i713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i712_3_lut (.I0(ram_s_3_3), .I1(register_vector[11]), .I2(n254), 
            .I3(GND_net), .O(n960));   // src/ram.vhd(56[12:17])
    defparam i712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i711_3_lut (.I0(ram_s_3_4), .I1(sx[4]), .I2(n254), .I3(GND_net), 
            .O(n959));   // src/ram.vhd(56[12:17])
    defparam i711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i710_3_lut (.I0(ram_s_3_5), .I1(sx[5]), .I2(n254), .I3(GND_net), 
            .O(n958));   // src/ram.vhd(56[12:17])
    defparam i710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i709_3_lut (.I0(ram_s_14_7), .I1(sx[7]), .I2(n243), .I3(GND_net), 
            .O(n957));   // src/ram.vhd(56[12:17])
    defparam i709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i704_3_lut (.I0(ram_s_3_6), .I1(sx[6]), .I2(n254), .I3(GND_net), 
            .O(n952));   // src/ram.vhd(56[12:17])
    defparam i704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i702_3_lut (.I0(ram_s_3_7), .I1(sx[7]), .I2(n254), .I3(GND_net), 
            .O(n950));   // src/ram.vhd(56[12:17])
    defparam i702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i698_3_lut (.I0(ram_s_4_0), .I1(register_vector[8]), .I2(n253), 
            .I3(GND_net), .O(n946));   // src/ram.vhd(56[12:17])
    defparam i698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i696_3_lut (.I0(ram_s_4_1), .I1(register_vector[9]), .I2(n253), 
            .I3(GND_net), .O(n944));   // src/ram.vhd(56[12:17])
    defparam i696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i693_3_lut (.I0(ram_s_4_2), .I1(register_vector[10]), .I2(n253), 
            .I3(GND_net), .O(n941));   // src/ram.vhd(56[12:17])
    defparam i693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i692_3_lut (.I0(ram_s_5_2), .I1(register_vector[10]), .I2(n252), 
            .I3(GND_net), .O(n940));   // src/ram.vhd(56[12:17])
    defparam i692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i691_3_lut (.I0(ram_s_5_3), .I1(register_vector[11]), .I2(n252), 
            .I3(GND_net), .O(n939));   // src/ram.vhd(56[12:17])
    defparam i691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i687_3_lut (.I0(ram_s_5_5), .I1(sx[5]), .I2(n252), .I3(GND_net), 
            .O(n935));   // src/ram.vhd(56[12:17])
    defparam i687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i686_3_lut (.I0(ram_s_6_0), .I1(register_vector[8]), .I2(n251), 
            .I3(GND_net), .O(n934));   // src/ram.vhd(56[12:17])
    defparam i686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i685_3_lut (.I0(ram_s_6_1), .I1(register_vector[9]), .I2(n251), 
            .I3(GND_net), .O(n933));   // src/ram.vhd(56[12:17])
    defparam i685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i684_3_lut (.I0(ram_s_6_2), .I1(register_vector[10]), .I2(n251), 
            .I3(GND_net), .O(n932));   // src/ram.vhd(56[12:17])
    defparam i684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i683_3_lut (.I0(ram_s_5_6), .I1(sx[6]), .I2(n252), .I3(GND_net), 
            .O(n931));   // src/ram.vhd(56[12:17])
    defparam i683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i682_3_lut (.I0(ram_s_5_7), .I1(sx[7]), .I2(n252), .I3(GND_net), 
            .O(n930));   // src/ram.vhd(56[12:17])
    defparam i682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i679_3_lut (.I0(ram_s_4_3), .I1(register_vector[11]), .I2(n253), 
            .I3(GND_net), .O(n927));   // src/ram.vhd(56[12:17])
    defparam i679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i678_3_lut (.I0(ram_s_13_5), .I1(sx[5]), .I2(n244), .I3(GND_net), 
            .O(n926));   // src/ram.vhd(56[12:17])
    defparam i678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i677_3_lut (.I0(ram_s_13_3), .I1(register_vector[11]), .I2(n244), 
            .I3(GND_net), .O(n925));   // src/ram.vhd(56[12:17])
    defparam i677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i676_3_lut (.I0(ram_s_13_4), .I1(sx[4]), .I2(n244), .I3(GND_net), 
            .O(n924));   // src/ram.vhd(56[12:17])
    defparam i676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i675_3_lut (.I0(ram_s_13_6), .I1(sx[6]), .I2(n244), .I3(GND_net), 
            .O(n923));   // src/ram.vhd(56[12:17])
    defparam i675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i690_4_lut_4_lut (.I0(internal_reset), .I1(address[0]), .I2(pc_value[0]), 
            .I3(t_state[1]), .O(n938));   // src/program_counter.vhd(55[9] 61[16])
    defparam i690_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i670_3_lut (.I0(ram_s_13_7), .I1(sx[7]), .I2(n244), .I3(GND_net), 
            .O(n918));   // src/ram.vhd(56[12:17])
    defparam i670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i669_3_lut (.I0(ram_s_14_0), .I1(register_vector[8]), .I2(n243), 
            .I3(GND_net), .O(n917));   // src/ram.vhd(56[12:17])
    defparam i669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i668_3_lut (.I0(ram_s_14_1), .I1(register_vector[9]), .I2(n243), 
            .I3(GND_net), .O(n916));   // src/ram.vhd(56[12:17])
    defparam i668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i663_3_lut (.I0(ram_s_13_2), .I1(register_vector[10]), .I2(n244), 
            .I3(GND_net), .O(n911));   // src/ram.vhd(56[12:17])
    defparam i663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i661_3_lut (.I0(ram_s_11_0), .I1(register_vector[8]), .I2(n246), 
            .I3(GND_net), .O(n909));   // src/ram.vhd(56[12:17])
    defparam i661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i660_3_lut (.I0(ram_s_14_3), .I1(register_vector[11]), .I2(n243), 
            .I3(GND_net), .O(n908));   // src/ram.vhd(56[12:17])
    defparam i660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i659_3_lut (.I0(ram_s_13_1), .I1(register_vector[9]), .I2(n244), 
            .I3(GND_net), .O(n907));   // src/ram.vhd(56[12:17])
    defparam i659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i658_3_lut (.I0(ram_s_14_2), .I1(register_vector[10]), .I2(n243), 
            .I3(GND_net), .O(n906));   // src/ram.vhd(56[12:17])
    defparam i658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i656_3_lut (.I0(ram_s_13_0), .I1(register_vector[8]), .I2(n244), 
            .I3(GND_net), .O(n904));   // src/ram.vhd(56[12:17])
    defparam i656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i653_3_lut (.I0(ram_s_5_4), .I1(sx[4]), .I2(n252), .I3(GND_net), 
            .O(n901));   // src/ram.vhd(56[12:17])
    defparam i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i651_3_lut (.I0(ram_s_14_6), .I1(sx[6]), .I2(n243), .I3(GND_net), 
            .O(n899));   // src/ram.vhd(56[12:17])
    defparam i651_3_lut.LUT_INIT = 16'hcaca;
    program_memory test_program (.wea({GND_net}), .VCC_net(VCC_net), .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), 
            .bram_enable(bram_enable), .\address[10] (address[10]), .\address[9] (address[9]), 
            .\address[8] (address[8]), .\address[7] (address[7]), .\address[6] (address[6]), 
            .\address[5] (address[5]), .\address[4] (address[4]), .\address[3] (address[3]), 
            .\address[2] (address[2]), .\address[1] (address[1]), .\address[0] (address[0]), 
            .instruction({instruction}));   // src/top.vhd(87[20:34])
    
endmodule
//
// Verilog Description of module zipi8
//

module zipi8 (CLK_3P3_MHZ_c, instruction, wea, \sx[7] , \sx[6] , \sx[5] , 
            \sx[4] , \register_vector[11] , \register_vector[10] , \register_vector[9] , 
            \register_vector[8] , n8580, bram_enable, \t_state[1] , 
            internal_reset, BTN1_c, special_bit, address, VCC_net, 
            ram_s_70_3, ram_s_71_3, ram_s_69_3, ram_s_68_3, ram_s_34_7, 
            ram_s_35_7, ram_s_33_7, ram_s_32_7, ram_s_11_6, ram_s_8_6, 
            ram_s_62_4, ram_s_63_4, ram_s_2_7, ram_s_3_7, ram_s_1_7, 
            ram_s_0_7, ram_s_66_4, ram_s_67_4, ram_s_65_4, ram_s_64_4, 
            ram_s_142_3, ram_s_141_3, ram_s_140_3, ram_s_209_3, ram_s_130_0, 
            ram_s_131_0, ram_s_129_0, ram_s_128_0, ram_s_70_4, ram_s_71_4, 
            ram_s_69_4, ram_s_68_4, ram_s_171_5, ram_s_168_5, ram_s_14_6, 
            ram_s_13_6, ram_s_12_6, ram_s_202_1, ram_s_203_1, ram_s_6_5, 
            ram_s_7_5, ram_s_14_5, ram_s_5_5, ram_s_4_5, ram_s_13_5, 
            ram_s_12_5, ram_s_43_2, ram_s_2_0, ram_s_3_0, ram_s_2_1, 
            ram_s_3_1, ram_s_1_0, ram_s_0_0, ram_s_66_0, ram_s_67_0, 
            ram_s_34_1, ram_s_35_1, ram_s_33_1, ram_s_32_1, ram_s_201_1, 
            ram_s_200_1, ram_s_1_1, ram_s_0_1, ram_s_65_0, ram_s_64_0, 
            ram_s_11_2, ram_s_8_2, ram_s_38_0, ram_s_39_0, ram_s_40_2, 
            ram_s_74_7, ram_s_75_7, ram_s_73_7, ram_s_72_7, ram_s_130_7, 
            ram_s_131_7, ram_s_129_7, ram_s_128_7, ram_s_37_0, ram_s_36_0, 
            ram_s_142_5, ram_s_141_5, ram_s_140_5, ram_s_62_0, ram_s_63_0, 
            ram_s_194_1, ram_s_195_1, ram_s_193_1, ram_s_192_1, ram_s_74_4, 
            ram_s_75_4, ram_s_73_4, ram_s_72_4, ram_s_43_7, ram_s_40_7, 
            ram_s_74_2, ram_s_75_2, ram_s_73_2, ram_s_72_2, ram_s_186_3, 
            ram_s_185_3, ram_s_190_2, ram_s_191_2, ram_s_43_1, ram_s_40_1, 
            ram_s_6_7, ram_s_7_7, ram_s_134_0, ram_s_135_0, ram_s_5_7, 
            ram_s_4_7, ram_s_133_0, ram_s_132_0, ram_s_34_2, ram_s_35_2, 
            ram_s_58_5, ram_s_58_0, ram_s_57_0, ram_s_139_0, ram_s_136_0, 
            ram_s_190_5, ram_s_191_5, ram_s_57_5, ram_s_33_2, ram_s_32_2, 
            ram_s_142_7, ram_s_141_7, ram_s_140_7, ram_s_81_5, ram_s_190_1, 
            ram_s_191_1, ram_s_139_1, ram_s_136_1, ram_s_38_7, ram_s_39_7, 
            ram_s_37_7, ram_s_36_7, n893, ram_s_14_4, ram_s_190_7, 
            ram_s_191_7, ram_s_47_2, ram_s_45_2, ram_s_44_2, ram_s_134_5, 
            ram_s_135_5, ram_s_133_5, ram_s_132_5, n2567, ram_s_209_7, 
            n2566, ram_s_209_6, n2565, ram_s_209_5, n2564, ram_s_209_4, 
            n2563, n2562, ram_s_209_2, n2561, ram_s_209_1, n2560, 
            ram_s_209_0, n2519, ram_s_203_7, n2518, ram_s_203_6, n2517, 
            ram_s_203_5, n2516, ram_s_203_4, n2515, ram_s_203_3, n2514, 
            ram_s_203_2, n2513, n2512, ram_s_203_0, n2511, ram_s_202_7, 
            n2510, ram_s_202_6, n2509, ram_s_202_5, n2508, ram_s_202_4, 
            n2507, ram_s_202_3, n2506, ram_s_202_2, n2505, n2504, 
            ram_s_202_0, n2503, ram_s_201_7, n2502, ram_s_201_6, n2501, 
            ram_s_201_5, n2500, ram_s_201_4, n2499, ram_s_201_3, n2498, 
            ram_s_201_2, n2497, n2496, ram_s_201_0, n2495, ram_s_200_7, 
            n2494, ram_s_200_6, n2493, ram_s_200_5, n2492, ram_s_200_4, 
            n2491, ram_s_200_3, n2490, ram_s_200_2, n2489, n2488, 
            ram_s_200_0, n2487, ram_s_199_7, n2486, ram_s_199_6, n2485, 
            ram_s_199_5, n2484, ram_s_199_4, n2483, ram_s_199_3, n2482, 
            ram_s_199_2, n2481, ram_s_199_1, n2480, ram_s_199_0, n2479, 
            ram_s_198_7, n2478, ram_s_198_6, n2477, ram_s_198_5, n2476, 
            ram_s_198_4, n2475, ram_s_198_3, n2474, ram_s_198_2, n2473, 
            ram_s_198_1, n2472, ram_s_198_0, n2471, ram_s_197_7, n2470, 
            ram_s_197_6, n2469, ram_s_197_5, n2468, ram_s_197_4, n2467, 
            ram_s_197_3, n2466, ram_s_197_2, n2465, ram_s_197_1, n2464, 
            ram_s_197_0, n2463, ram_s_196_7, n2462, ram_s_196_6, n2461, 
            ram_s_196_5, n2460, ram_s_196_4, n2459, ram_s_196_3, n2458, 
            ram_s_196_2, n2457, ram_s_196_1, n2456, ram_s_196_0, n2455, 
            ram_s_195_7, n2454, ram_s_195_6, n2453, ram_s_195_5, n2452, 
            ram_s_195_4, n2451, ram_s_195_3, n2450, ram_s_195_2, n2449, 
            n2448, ram_s_195_0, n2447, ram_s_194_7, n2446, ram_s_194_6, 
            n2445, ram_s_194_5, n2444, ram_s_194_4, n2443, ram_s_194_3, 
            n2442, ram_s_194_2, n2441, n2440, ram_s_194_0, n2439, 
            ram_s_193_7, n2438, ram_s_193_6, n2437, ram_s_193_5, n2436, 
            ram_s_193_4, n2435, ram_s_193_3, n2434, ram_s_193_2, n2433, 
            n2432, ram_s_193_0, n2431, ram_s_192_7, n2430, ram_s_192_6, 
            n2429, ram_s_192_5, n2428, ram_s_192_4, n2427, ram_s_192_3, 
            n2426, ram_s_192_2, n2425, n2424, ram_s_192_0, n2423, 
            n2422, ram_s_191_6, n2421, n2420, ram_s_191_4, n2419, 
            ram_s_191_3, n2418, n2417, n2416, ram_s_191_0, n2415, 
            n2414, ram_s_190_6, n2413, n2412, ram_s_190_4, n2411, 
            ram_s_190_3, n2410, n2409, n2408, ram_s_190_0, n2383, 
            ram_s_186_7, n2382, ram_s_186_6, n2381, ram_s_186_5, n2380, 
            ram_s_186_4, n2379, n2378, ram_s_186_2, n2377, ram_s_186_1, 
            n2376, ram_s_186_0, n2375, ram_s_185_7, n2374, ram_s_185_6, 
            n2373, ram_s_185_5, n2372, ram_s_185_4, n2371, n2370, 
            ram_s_185_2, n2369, ram_s_185_1, n2368, ram_s_185_0, n2295, 
            ram_s_175_7, n2294, ram_s_175_6, n2293, ram_s_175_5, n2292, 
            ram_s_175_4, n2291, ram_s_175_3, n2290, ram_s_175_2, n2289, 
            ram_s_175_1, n2288, ram_s_175_0, n2279, ram_s_173_7, n2278, 
            ram_s_173_6, n2277, ram_s_173_5, n2276, ram_s_173_4, n2275, 
            ram_s_173_3, n2274, ram_s_173_2, n2273, ram_s_173_1, n2272, 
            ram_s_173_0, n2271, ram_s_172_7, n2270, ram_s_172_6, n2269, 
            ram_s_172_5, n2268, ram_s_172_4, n2267, ram_s_172_3, n2266, 
            ram_s_172_2, n2265, ram_s_172_1, n2264, ram_s_172_0, n2263, 
            ram_s_171_7, n2262, ram_s_171_6, n2261, n2260, ram_s_171_4, 
            n2259, ram_s_171_3, n2258, ram_s_171_2, n2257, ram_s_171_1, 
            n2256, ram_s_171_0, n2239, ram_s_168_7, n2238, ram_s_168_6, 
            n2237, n2236, ram_s_168_4, n2235, ram_s_168_3, n2234, 
            ram_s_168_2, n2233, ram_s_168_1, n2232, ram_s_168_0, n2231, 
            ram_s_167_7, n2230, ram_s_167_6, n2229, ram_s_167_5, n2228, 
            ram_s_167_4, n2227, ram_s_167_3, n2226, ram_s_167_2, n2225, 
            ram_s_167_1, n2224, ram_s_167_0, n2223, ram_s_166_7, n2222, 
            ram_s_166_6, n2221, ram_s_166_5, n2220, ram_s_166_4, n2219, 
            ram_s_166_3, n2218, ram_s_166_2, n2217, ram_s_166_1, n2216, 
            ram_s_166_0, n2215, ram_s_165_7, n2214, ram_s_165_6, n2213, 
            ram_s_165_5, n2212, ram_s_165_4, n2211, ram_s_165_3, n2210, 
            ram_s_165_2, n2209, ram_s_165_1, n2208, ram_s_165_0, n2207, 
            ram_s_164_7, n2206, ram_s_164_6, n2205, ram_s_164_5, n2204, 
            ram_s_164_4, n2203, ram_s_164_3, n2202, ram_s_164_2, n2201, 
            ram_s_164_1, n2200, ram_s_164_0, n2199, ram_s_163_7, n2198, 
            ram_s_163_6, n2197, ram_s_163_5, n2196, ram_s_163_4, n2195, 
            ram_s_163_3, n2194, ram_s_163_2, n2193, ram_s_163_1, n2192, 
            ram_s_163_0, n2191, ram_s_162_7, n2190, ram_s_162_6, n2189, 
            ram_s_162_5, n2188, ram_s_162_4, n2187, ram_s_162_3, n2186, 
            ram_s_162_2, n2185, ram_s_162_1, n2184, ram_s_162_0, n2183, 
            ram_s_161_7, n2182, ram_s_161_6, n2181, ram_s_161_5, n2180, 
            ram_s_161_4, n2179, ram_s_161_3, n2178, ram_s_161_2, n2177, 
            ram_s_161_1, n2176, ram_s_161_0, n2175, ram_s_160_7, n2174, 
            ram_s_160_6, n2173, ram_s_160_5, n2172, ram_s_160_4, n2171, 
            ram_s_160_3, n2170, ram_s_160_2, n2169, ram_s_160_1, n2168, 
            ram_s_160_0, n2031, n2030, ram_s_142_6, n2029, n2028, 
            ram_s_142_4, n2027, n2026, ram_s_142_2, n2025, ram_s_142_1, 
            n2024, ram_s_142_0, n2023, n2022, ram_s_141_6, n2021, 
            n2020, ram_s_141_4, n2019, n2018, ram_s_141_2, n2017, 
            ram_s_141_1, n2016, ram_s_141_0, n2015, n2014, ram_s_140_6, 
            n2013, n2012, ram_s_140_4, n2011, n2010, ram_s_140_2, 
            n2009, ram_s_140_1, n2008, ram_s_140_0, n2007, ram_s_139_7, 
            n2006, ram_s_139_6, n2005, ram_s_139_5, n2004, ram_s_139_4, 
            n2003, ram_s_139_3, n2002, ram_s_139_2, n2001, n2000, 
            n1983, ram_s_136_7, n1982, ram_s_136_6, n1981, ram_s_136_5, 
            n1980, ram_s_136_4, n1979, ram_s_136_3, n1978, ram_s_136_2, 
            n1977, n1976, n1975, ram_s_135_7, n1974, ram_s_135_6, 
            n1973, n1972, ram_s_135_4, n1971, ram_s_135_3, n1970, 
            ram_s_135_2, n1969, ram_s_135_1, n1968, n1967, ram_s_134_7, 
            n1966, ram_s_134_6, n1965, n1964, ram_s_134_4, n1963, 
            ram_s_134_3, n1962, ram_s_134_2, n1961, ram_s_134_1, n1960, 
            n1959, ram_s_133_7, n1958, ram_s_133_6, n1957, n1956, 
            ram_s_133_4, n1955, ram_s_133_3, n1954, ram_s_133_2, n1953, 
            ram_s_133_1, n1952, n1951, ram_s_132_7, n1950, ram_s_132_6, 
            n1949, n1948, ram_s_132_4, n1947, ram_s_132_3, n1946, 
            ram_s_132_2, n1945, ram_s_132_1, n1944, n1943, n1942, 
            ram_s_131_6, n1941, ram_s_131_5, n1940, ram_s_131_4, n1939, 
            ram_s_131_3, n1938, ram_s_131_2, n1937, ram_s_131_1, n1936, 
            n1935, n1934, ram_s_130_6, n1933, ram_s_130_5, n1932, 
            ram_s_130_4, n1931, ram_s_130_3, n1930, ram_s_130_2, n1929, 
            ram_s_130_1, n1928, n1927, n1926, ram_s_129_6, n1925, 
            ram_s_129_5, n1924, ram_s_129_4, n1923, ram_s_129_3, n1922, 
            ram_s_129_2, n1921, ram_s_129_1, n1920, n1919, n1918, 
            ram_s_128_6, n1917, ram_s_128_5, n1916, ram_s_128_4, n1915, 
            ram_s_128_3, n1914, ram_s_128_2, n1913, ram_s_128_1, n1912, 
            n1543, ram_s_81_7, n1542, ram_s_81_6, n1541, n1540, 
            ram_s_81_4, n1539, ram_s_81_3, n1538, ram_s_81_2, n1537, 
            ram_s_81_1, n1536, ram_s_81_0, n1495, n1494, ram_s_75_6, 
            n1493, ram_s_75_5, n1492, n1491, ram_s_75_3, n1490, 
            n1489, ram_s_75_1, n1488, ram_s_75_0, n1487, n1486, 
            ram_s_74_6, n1485, ram_s_74_5, n1484, n1483, ram_s_74_3, 
            n1482, n1481, ram_s_74_1, n1480, ram_s_74_0, n1479, 
            n1478, ram_s_73_6, n1477, ram_s_73_5, n1476, n1475, 
            ram_s_73_3, n1474, n1473, ram_s_73_1, n1472, ram_s_73_0, 
            n1471, n1470, ram_s_72_6, n1469, ram_s_72_5, n1468, 
            n1467, ram_s_72_3, n1466, n1465, ram_s_72_1, n1464, 
            ram_s_72_0, n1463, ram_s_71_7, n1462, ram_s_71_6, n1461, 
            ram_s_71_5, n1460, n1459, n1458, ram_s_71_2, n1457, 
            ram_s_71_1, n1456, ram_s_71_0, n1455, ram_s_70_7, n1454, 
            ram_s_70_6, n1453, ram_s_70_5, n1452, n1451, n1450, 
            ram_s_70_2, n1449, ram_s_70_1, n1448, ram_s_70_0, n1447, 
            ram_s_69_7, n1446, ram_s_69_6, n1445, ram_s_69_5, n1444, 
            n1443, n1442, ram_s_69_2, n1441, ram_s_69_1, n1440, 
            ram_s_69_0, n1439, ram_s_68_7, n1438, ram_s_68_6, n1437, 
            ram_s_68_5, n1436, n1435, n1434, ram_s_68_2, n1433, 
            ram_s_68_1, n1432, ram_s_68_0, n1431, ram_s_67_7, n1430, 
            ram_s_67_6, n1429, ram_s_67_5, n1428, n1427, ram_s_67_3, 
            n1426, ram_s_67_2, n1425, ram_s_67_1, n1424, n1423, 
            ram_s_66_7, n1422, ram_s_66_6, n1421, ram_s_66_5, n1420, 
            n1419, ram_s_66_3, n1418, ram_s_66_2, n1417, ram_s_66_1, 
            n1416, n1415, ram_s_65_7, n1414, ram_s_65_6, n1413, 
            ram_s_65_5, n1412, n1411, ram_s_65_3, n1410, ram_s_65_2, 
            n1409, ram_s_65_1, n1408, n1407, ram_s_64_7, n1406, 
            ram_s_64_6, n1405, ram_s_64_5, n1404, n1403, ram_s_64_3, 
            n1402, ram_s_64_2, n1401, ram_s_64_1, n1400, n1399, 
            ram_s_63_7, n1398, ram_s_63_6, n1397, ram_s_63_5, n1396, 
            n1395, ram_s_63_3, n1394, ram_s_63_2, n1393, ram_s_63_1, 
            n1392, n1391, ram_s_62_7, n1390, ram_s_62_6, n1389, 
            ram_s_62_5, n1388, n1387, ram_s_62_3, n1386, ram_s_62_2, 
            n1385, ram_s_62_1, n1384, n1359, ram_s_58_7, n1358, 
            ram_s_58_6, n1357, n1356, ram_s_58_4, n1355, ram_s_58_3, 
            n1354, ram_s_58_2, n1353, ram_s_58_1, n1352, n1351, 
            ram_s_57_7, n1350, ram_s_57_6, n1349, n1348, ram_s_57_4, 
            n1347, ram_s_57_3, n1346, ram_s_57_2, n1345, ram_s_57_1, 
            n1344, n1271, ram_s_47_7, n1270, ram_s_47_6, n1269, 
            ram_s_47_5, n1268, ram_s_47_4, n1267, ram_s_47_3, n1266, 
            n1265, ram_s_47_1, n1264, ram_s_47_0, n1255, ram_s_45_7, 
            n1254, ram_s_45_6, n1253, ram_s_45_5, n1252, ram_s_45_4, 
            n1251, ram_s_45_3, n1250, n1249, ram_s_45_1, n1248, 
            ram_s_45_0, n1247, ram_s_44_7, n1246, ram_s_44_6, n1245, 
            ram_s_44_5, n1244, ram_s_44_4, n1243, ram_s_44_3, n1242, 
            n1241, ram_s_44_1, n1240, ram_s_44_0, n1239, n1238, 
            ram_s_43_6, n1237, ram_s_43_5, n1236, ram_s_43_4, n1235, 
            ram_s_43_3, n1234, n1233, n1232, ram_s_43_0, n1215, 
            n1214, ram_s_40_6, n1213, ram_s_40_5, n1212, ram_s_40_4, 
            n1211, ram_s_40_3, n1210, n1209, n1208, ram_s_40_0, 
            n1207, n1206, ram_s_39_6, n1205, ram_s_39_5, n1204, 
            ram_s_39_4, n1203, ram_s_39_3, n1202, ram_s_39_2, n1201, 
            ram_s_39_1, n1200, n1199, n1198, ram_s_38_6, n1197, 
            ram_s_38_5, n1196, ram_s_38_4, n1195, ram_s_38_3, n1194, 
            ram_s_38_2, n1193, ram_s_38_1, n1192, n1191, n1190, 
            ram_s_37_6, n1189, ram_s_37_5, n1188, ram_s_37_4, n1187, 
            ram_s_37_3, n1186, ram_s_37_2, n1185, ram_s_37_1, n1184, 
            n1183, n1182, ram_s_36_6, n1181, ram_s_36_5, n1180, 
            ram_s_36_4, n1179, ram_s_36_3, n1178, ram_s_36_2, n1177, 
            ram_s_36_1, n1176, n1175, n1174, ram_s_35_6, n1173, 
            ram_s_35_5, n1172, ram_s_35_4, n1171, ram_s_35_3, n1170, 
            n1169, n1168, ram_s_35_0, n1167, n1166, ram_s_34_6, 
            n1165, ram_s_34_5, n1164, ram_s_34_4, n1163, ram_s_34_3, 
            n1162, n1161, n1160, ram_s_34_0, n1159, n1158, ram_s_33_6, 
            n1157, ram_s_33_5, n1156, ram_s_33_4, n1155, ram_s_33_3, 
            n1154, n1153, n1152, ram_s_33_0, n1151, n1150, ram_s_32_6, 
            n1149, ram_s_32_5, n1148, ram_s_32_4, n1147, ram_s_32_3, 
            n1146, n1145, n1144, ram_s_32_0, n1051, n1047, n1046, 
            n1045, ram_s_0_2, n1044, ram_s_12_3, n1043, n1042, ram_s_11_1, 
            n1041, n1040, ram_s_12_1, n1038, ram_s_11_4, n182, n1037, 
            ram_s_12_4, n54, n1036, ram_s_11_7, n183, n1035, n55, 
            n1034, ram_s_12_7, n184, n1033, ram_s_12_2, n56, n1032, 
            ram_s_11_5, n185, n1031, n57, n1030, ram_s_12_0, n186, 
            n1029, ram_s_11_3, n58, n187, n59, n188, n60, n189, 
            n61, n190, n62, n191, n63, n192, n1017, ram_s_0_3, 
            n64, n1016, ram_s_0_4, n193, n1015, ram_s_0_5, n65, 
            n1014, ram_s_0_6, n194, n1013, n66, n1012, n195, n1011, 
            n67, n1010, ram_s_1_2, n1009, ram_s_1_3, n1008, ram_s_1_4, 
            n1007, ram_s_1_5, n1006, ram_s_4_4, n1005, n1004, n1003, 
            ram_s_5_0, n1002, ram_s_4_6, n1001, ram_s_5_1, n998, 
            ram_s_8_5, n997, n996, n995, ram_s_7_4, n994, ram_s_7_1, 
            n993, ram_s_6_6, n992, ram_s_6_3, n989, n988, ram_s_8_3, 
            n987, ram_s_8_0, n986, n199, n985, ram_s_7_2, n71, 
            n984, n200, n983, ram_s_6_4, n72, n980, ram_s_8_7, 
            n979, ram_s_8_4, n978, ram_s_8_1, n977, ram_s_7_6, n976, 
            ram_s_7_3, n975, ram_s_7_0, n974, n973, ram_s_1_6, n972, 
            n971, n970, n969, ram_s_2_2, n968, ram_s_2_3, n967, 
            ram_s_2_4, n966, ram_s_2_5, n965, ram_s_2_6, n964, n963, 
            n962, n961, ram_s_3_2, n960, ram_s_3_3, n959, ram_s_3_4, 
            n958, ram_s_3_5, n957, ram_s_14_7, n952, ram_s_3_6, 
            n950, n946, ram_s_4_0, n944, ram_s_4_1, n941, ram_s_4_2, 
            n940, ram_s_5_2, n939, ram_s_5_3, n935, n934, ram_s_6_0, 
            n933, ram_s_6_1, n932, ram_s_6_2, n931, ram_s_5_6, n930, 
            n927, ram_s_4_3, n926, n925, ram_s_13_3, n924, ram_s_13_4, 
            n923, n210, n82, n212, n84, n213, n85, n214, n86, 
            n217, n89, n218, n90, n219, n91, n220, n92, n221, 
            n93, n222, n94, n223, n95, n224, n96, n225, n97, 
            n918, ram_s_13_7, n917, ram_s_14_0, n916, ram_s_14_1, 
            n244, n116, n115, n243, n245, n117, n246, n118, 
            n48, n176, n249, n121, n250, n122, n251, n123, n252, 
            n124, n253, n125, n254, n126, n255, n127, n256, 
            n128, n257, n129, ram_s_14_2, ram_s_13_2, ram_s_11_0, 
            n911, n909, n908, ram_s_14_3, n907, ram_s_13_1, n906, 
            n904, ram_s_13_0, n901, ram_s_5_4, n899, LED1_c_0, n765, 
            n938, \pc_value[0] );
    input CLK_3P3_MHZ_c;
    input [17:0]instruction;
    input [0:0]wea;
    output \sx[7] ;
    output \sx[6] ;
    output \sx[5] ;
    output \sx[4] ;
    output \register_vector[11] ;
    output \register_vector[10] ;
    output \register_vector[9] ;
    output \register_vector[8] ;
    input n8580;
    output bram_enable;
    output \t_state[1] ;
    output internal_reset;
    input BTN1_c;
    output special_bit;
    output [11:0]address;
    input VCC_net;
    output ram_s_70_3;
    output ram_s_71_3;
    output ram_s_69_3;
    output ram_s_68_3;
    output ram_s_34_7;
    output ram_s_35_7;
    output ram_s_33_7;
    output ram_s_32_7;
    output ram_s_11_6;
    output ram_s_8_6;
    output ram_s_62_4;
    output ram_s_63_4;
    output ram_s_2_7;
    output ram_s_3_7;
    output ram_s_1_7;
    output ram_s_0_7;
    output ram_s_66_4;
    output ram_s_67_4;
    output ram_s_65_4;
    output ram_s_64_4;
    output ram_s_142_3;
    output ram_s_141_3;
    output ram_s_140_3;
    output ram_s_209_3;
    output ram_s_130_0;
    output ram_s_131_0;
    output ram_s_129_0;
    output ram_s_128_0;
    output ram_s_70_4;
    output ram_s_71_4;
    output ram_s_69_4;
    output ram_s_68_4;
    output ram_s_171_5;
    output ram_s_168_5;
    output ram_s_14_6;
    output ram_s_13_6;
    output ram_s_12_6;
    output ram_s_202_1;
    output ram_s_203_1;
    output ram_s_6_5;
    output ram_s_7_5;
    output ram_s_14_5;
    output ram_s_5_5;
    output ram_s_4_5;
    output ram_s_13_5;
    output ram_s_12_5;
    output ram_s_43_2;
    output ram_s_2_0;
    output ram_s_3_0;
    output ram_s_2_1;
    output ram_s_3_1;
    output ram_s_1_0;
    output ram_s_0_0;
    output ram_s_66_0;
    output ram_s_67_0;
    output ram_s_34_1;
    output ram_s_35_1;
    output ram_s_33_1;
    output ram_s_32_1;
    output ram_s_201_1;
    output ram_s_200_1;
    output ram_s_1_1;
    output ram_s_0_1;
    output ram_s_65_0;
    output ram_s_64_0;
    output ram_s_11_2;
    output ram_s_8_2;
    output ram_s_38_0;
    output ram_s_39_0;
    output ram_s_40_2;
    output ram_s_74_7;
    output ram_s_75_7;
    output ram_s_73_7;
    output ram_s_72_7;
    output ram_s_130_7;
    output ram_s_131_7;
    output ram_s_129_7;
    output ram_s_128_7;
    output ram_s_37_0;
    output ram_s_36_0;
    output ram_s_142_5;
    output ram_s_141_5;
    output ram_s_140_5;
    output ram_s_62_0;
    output ram_s_63_0;
    output ram_s_194_1;
    output ram_s_195_1;
    output ram_s_193_1;
    output ram_s_192_1;
    output ram_s_74_4;
    output ram_s_75_4;
    output ram_s_73_4;
    output ram_s_72_4;
    output ram_s_43_7;
    output ram_s_40_7;
    output ram_s_74_2;
    output ram_s_75_2;
    output ram_s_73_2;
    output ram_s_72_2;
    output ram_s_186_3;
    output ram_s_185_3;
    output ram_s_190_2;
    output ram_s_191_2;
    output ram_s_43_1;
    output ram_s_40_1;
    output ram_s_6_7;
    output ram_s_7_7;
    output ram_s_134_0;
    output ram_s_135_0;
    output ram_s_5_7;
    output ram_s_4_7;
    output ram_s_133_0;
    output ram_s_132_0;
    output ram_s_34_2;
    output ram_s_35_2;
    output ram_s_58_5;
    output ram_s_58_0;
    output ram_s_57_0;
    output ram_s_139_0;
    output ram_s_136_0;
    output ram_s_190_5;
    output ram_s_191_5;
    output ram_s_57_5;
    output ram_s_33_2;
    output ram_s_32_2;
    output ram_s_142_7;
    output ram_s_141_7;
    output ram_s_140_7;
    output ram_s_81_5;
    output ram_s_190_1;
    output ram_s_191_1;
    output ram_s_139_1;
    output ram_s_136_1;
    output ram_s_38_7;
    output ram_s_39_7;
    output ram_s_37_7;
    output ram_s_36_7;
    input n893;
    output ram_s_14_4;
    output ram_s_190_7;
    output ram_s_191_7;
    output ram_s_47_2;
    output ram_s_45_2;
    output ram_s_44_2;
    output ram_s_134_5;
    output ram_s_135_5;
    output ram_s_133_5;
    output ram_s_132_5;
    input n2567;
    output ram_s_209_7;
    input n2566;
    output ram_s_209_6;
    input n2565;
    output ram_s_209_5;
    input n2564;
    output ram_s_209_4;
    input n2563;
    input n2562;
    output ram_s_209_2;
    input n2561;
    output ram_s_209_1;
    input n2560;
    output ram_s_209_0;
    input n2519;
    output ram_s_203_7;
    input n2518;
    output ram_s_203_6;
    input n2517;
    output ram_s_203_5;
    input n2516;
    output ram_s_203_4;
    input n2515;
    output ram_s_203_3;
    input n2514;
    output ram_s_203_2;
    input n2513;
    input n2512;
    output ram_s_203_0;
    input n2511;
    output ram_s_202_7;
    input n2510;
    output ram_s_202_6;
    input n2509;
    output ram_s_202_5;
    input n2508;
    output ram_s_202_4;
    input n2507;
    output ram_s_202_3;
    input n2506;
    output ram_s_202_2;
    input n2505;
    input n2504;
    output ram_s_202_0;
    input n2503;
    output ram_s_201_7;
    input n2502;
    output ram_s_201_6;
    input n2501;
    output ram_s_201_5;
    input n2500;
    output ram_s_201_4;
    input n2499;
    output ram_s_201_3;
    input n2498;
    output ram_s_201_2;
    input n2497;
    input n2496;
    output ram_s_201_0;
    input n2495;
    output ram_s_200_7;
    input n2494;
    output ram_s_200_6;
    input n2493;
    output ram_s_200_5;
    input n2492;
    output ram_s_200_4;
    input n2491;
    output ram_s_200_3;
    input n2490;
    output ram_s_200_2;
    input n2489;
    input n2488;
    output ram_s_200_0;
    input n2487;
    output ram_s_199_7;
    input n2486;
    output ram_s_199_6;
    input n2485;
    output ram_s_199_5;
    input n2484;
    output ram_s_199_4;
    input n2483;
    output ram_s_199_3;
    input n2482;
    output ram_s_199_2;
    input n2481;
    output ram_s_199_1;
    input n2480;
    output ram_s_199_0;
    input n2479;
    output ram_s_198_7;
    input n2478;
    output ram_s_198_6;
    input n2477;
    output ram_s_198_5;
    input n2476;
    output ram_s_198_4;
    input n2475;
    output ram_s_198_3;
    input n2474;
    output ram_s_198_2;
    input n2473;
    output ram_s_198_1;
    input n2472;
    output ram_s_198_0;
    input n2471;
    output ram_s_197_7;
    input n2470;
    output ram_s_197_6;
    input n2469;
    output ram_s_197_5;
    input n2468;
    output ram_s_197_4;
    input n2467;
    output ram_s_197_3;
    input n2466;
    output ram_s_197_2;
    input n2465;
    output ram_s_197_1;
    input n2464;
    output ram_s_197_0;
    input n2463;
    output ram_s_196_7;
    input n2462;
    output ram_s_196_6;
    input n2461;
    output ram_s_196_5;
    input n2460;
    output ram_s_196_4;
    input n2459;
    output ram_s_196_3;
    input n2458;
    output ram_s_196_2;
    input n2457;
    output ram_s_196_1;
    input n2456;
    output ram_s_196_0;
    input n2455;
    output ram_s_195_7;
    input n2454;
    output ram_s_195_6;
    input n2453;
    output ram_s_195_5;
    input n2452;
    output ram_s_195_4;
    input n2451;
    output ram_s_195_3;
    input n2450;
    output ram_s_195_2;
    input n2449;
    input n2448;
    output ram_s_195_0;
    input n2447;
    output ram_s_194_7;
    input n2446;
    output ram_s_194_6;
    input n2445;
    output ram_s_194_5;
    input n2444;
    output ram_s_194_4;
    input n2443;
    output ram_s_194_3;
    input n2442;
    output ram_s_194_2;
    input n2441;
    input n2440;
    output ram_s_194_0;
    input n2439;
    output ram_s_193_7;
    input n2438;
    output ram_s_193_6;
    input n2437;
    output ram_s_193_5;
    input n2436;
    output ram_s_193_4;
    input n2435;
    output ram_s_193_3;
    input n2434;
    output ram_s_193_2;
    input n2433;
    input n2432;
    output ram_s_193_0;
    input n2431;
    output ram_s_192_7;
    input n2430;
    output ram_s_192_6;
    input n2429;
    output ram_s_192_5;
    input n2428;
    output ram_s_192_4;
    input n2427;
    output ram_s_192_3;
    input n2426;
    output ram_s_192_2;
    input n2425;
    input n2424;
    output ram_s_192_0;
    input n2423;
    input n2422;
    output ram_s_191_6;
    input n2421;
    input n2420;
    output ram_s_191_4;
    input n2419;
    output ram_s_191_3;
    input n2418;
    input n2417;
    input n2416;
    output ram_s_191_0;
    input n2415;
    input n2414;
    output ram_s_190_6;
    input n2413;
    input n2412;
    output ram_s_190_4;
    input n2411;
    output ram_s_190_3;
    input n2410;
    input n2409;
    input n2408;
    output ram_s_190_0;
    input n2383;
    output ram_s_186_7;
    input n2382;
    output ram_s_186_6;
    input n2381;
    output ram_s_186_5;
    input n2380;
    output ram_s_186_4;
    input n2379;
    input n2378;
    output ram_s_186_2;
    input n2377;
    output ram_s_186_1;
    input n2376;
    output ram_s_186_0;
    input n2375;
    output ram_s_185_7;
    input n2374;
    output ram_s_185_6;
    input n2373;
    output ram_s_185_5;
    input n2372;
    output ram_s_185_4;
    input n2371;
    input n2370;
    output ram_s_185_2;
    input n2369;
    output ram_s_185_1;
    input n2368;
    output ram_s_185_0;
    input n2295;
    output ram_s_175_7;
    input n2294;
    output ram_s_175_6;
    input n2293;
    output ram_s_175_5;
    input n2292;
    output ram_s_175_4;
    input n2291;
    output ram_s_175_3;
    input n2290;
    output ram_s_175_2;
    input n2289;
    output ram_s_175_1;
    input n2288;
    output ram_s_175_0;
    input n2279;
    output ram_s_173_7;
    input n2278;
    output ram_s_173_6;
    input n2277;
    output ram_s_173_5;
    input n2276;
    output ram_s_173_4;
    input n2275;
    output ram_s_173_3;
    input n2274;
    output ram_s_173_2;
    input n2273;
    output ram_s_173_1;
    input n2272;
    output ram_s_173_0;
    input n2271;
    output ram_s_172_7;
    input n2270;
    output ram_s_172_6;
    input n2269;
    output ram_s_172_5;
    input n2268;
    output ram_s_172_4;
    input n2267;
    output ram_s_172_3;
    input n2266;
    output ram_s_172_2;
    input n2265;
    output ram_s_172_1;
    input n2264;
    output ram_s_172_0;
    input n2263;
    output ram_s_171_7;
    input n2262;
    output ram_s_171_6;
    input n2261;
    input n2260;
    output ram_s_171_4;
    input n2259;
    output ram_s_171_3;
    input n2258;
    output ram_s_171_2;
    input n2257;
    output ram_s_171_1;
    input n2256;
    output ram_s_171_0;
    input n2239;
    output ram_s_168_7;
    input n2238;
    output ram_s_168_6;
    input n2237;
    input n2236;
    output ram_s_168_4;
    input n2235;
    output ram_s_168_3;
    input n2234;
    output ram_s_168_2;
    input n2233;
    output ram_s_168_1;
    input n2232;
    output ram_s_168_0;
    input n2231;
    output ram_s_167_7;
    input n2230;
    output ram_s_167_6;
    input n2229;
    output ram_s_167_5;
    input n2228;
    output ram_s_167_4;
    input n2227;
    output ram_s_167_3;
    input n2226;
    output ram_s_167_2;
    input n2225;
    output ram_s_167_1;
    input n2224;
    output ram_s_167_0;
    input n2223;
    output ram_s_166_7;
    input n2222;
    output ram_s_166_6;
    input n2221;
    output ram_s_166_5;
    input n2220;
    output ram_s_166_4;
    input n2219;
    output ram_s_166_3;
    input n2218;
    output ram_s_166_2;
    input n2217;
    output ram_s_166_1;
    input n2216;
    output ram_s_166_0;
    input n2215;
    output ram_s_165_7;
    input n2214;
    output ram_s_165_6;
    input n2213;
    output ram_s_165_5;
    input n2212;
    output ram_s_165_4;
    input n2211;
    output ram_s_165_3;
    input n2210;
    output ram_s_165_2;
    input n2209;
    output ram_s_165_1;
    input n2208;
    output ram_s_165_0;
    input n2207;
    output ram_s_164_7;
    input n2206;
    output ram_s_164_6;
    input n2205;
    output ram_s_164_5;
    input n2204;
    output ram_s_164_4;
    input n2203;
    output ram_s_164_3;
    input n2202;
    output ram_s_164_2;
    input n2201;
    output ram_s_164_1;
    input n2200;
    output ram_s_164_0;
    input n2199;
    output ram_s_163_7;
    input n2198;
    output ram_s_163_6;
    input n2197;
    output ram_s_163_5;
    input n2196;
    output ram_s_163_4;
    input n2195;
    output ram_s_163_3;
    input n2194;
    output ram_s_163_2;
    input n2193;
    output ram_s_163_1;
    input n2192;
    output ram_s_163_0;
    input n2191;
    output ram_s_162_7;
    input n2190;
    output ram_s_162_6;
    input n2189;
    output ram_s_162_5;
    input n2188;
    output ram_s_162_4;
    input n2187;
    output ram_s_162_3;
    input n2186;
    output ram_s_162_2;
    input n2185;
    output ram_s_162_1;
    input n2184;
    output ram_s_162_0;
    input n2183;
    output ram_s_161_7;
    input n2182;
    output ram_s_161_6;
    input n2181;
    output ram_s_161_5;
    input n2180;
    output ram_s_161_4;
    input n2179;
    output ram_s_161_3;
    input n2178;
    output ram_s_161_2;
    input n2177;
    output ram_s_161_1;
    input n2176;
    output ram_s_161_0;
    input n2175;
    output ram_s_160_7;
    input n2174;
    output ram_s_160_6;
    input n2173;
    output ram_s_160_5;
    input n2172;
    output ram_s_160_4;
    input n2171;
    output ram_s_160_3;
    input n2170;
    output ram_s_160_2;
    input n2169;
    output ram_s_160_1;
    input n2168;
    output ram_s_160_0;
    input n2031;
    input n2030;
    output ram_s_142_6;
    input n2029;
    input n2028;
    output ram_s_142_4;
    input n2027;
    input n2026;
    output ram_s_142_2;
    input n2025;
    output ram_s_142_1;
    input n2024;
    output ram_s_142_0;
    input n2023;
    input n2022;
    output ram_s_141_6;
    input n2021;
    input n2020;
    output ram_s_141_4;
    input n2019;
    input n2018;
    output ram_s_141_2;
    input n2017;
    output ram_s_141_1;
    input n2016;
    output ram_s_141_0;
    input n2015;
    input n2014;
    output ram_s_140_6;
    input n2013;
    input n2012;
    output ram_s_140_4;
    input n2011;
    input n2010;
    output ram_s_140_2;
    input n2009;
    output ram_s_140_1;
    input n2008;
    output ram_s_140_0;
    input n2007;
    output ram_s_139_7;
    input n2006;
    output ram_s_139_6;
    input n2005;
    output ram_s_139_5;
    input n2004;
    output ram_s_139_4;
    input n2003;
    output ram_s_139_3;
    input n2002;
    output ram_s_139_2;
    input n2001;
    input n2000;
    input n1983;
    output ram_s_136_7;
    input n1982;
    output ram_s_136_6;
    input n1981;
    output ram_s_136_5;
    input n1980;
    output ram_s_136_4;
    input n1979;
    output ram_s_136_3;
    input n1978;
    output ram_s_136_2;
    input n1977;
    input n1976;
    input n1975;
    output ram_s_135_7;
    input n1974;
    output ram_s_135_6;
    input n1973;
    input n1972;
    output ram_s_135_4;
    input n1971;
    output ram_s_135_3;
    input n1970;
    output ram_s_135_2;
    input n1969;
    output ram_s_135_1;
    input n1968;
    input n1967;
    output ram_s_134_7;
    input n1966;
    output ram_s_134_6;
    input n1965;
    input n1964;
    output ram_s_134_4;
    input n1963;
    output ram_s_134_3;
    input n1962;
    output ram_s_134_2;
    input n1961;
    output ram_s_134_1;
    input n1960;
    input n1959;
    output ram_s_133_7;
    input n1958;
    output ram_s_133_6;
    input n1957;
    input n1956;
    output ram_s_133_4;
    input n1955;
    output ram_s_133_3;
    input n1954;
    output ram_s_133_2;
    input n1953;
    output ram_s_133_1;
    input n1952;
    input n1951;
    output ram_s_132_7;
    input n1950;
    output ram_s_132_6;
    input n1949;
    input n1948;
    output ram_s_132_4;
    input n1947;
    output ram_s_132_3;
    input n1946;
    output ram_s_132_2;
    input n1945;
    output ram_s_132_1;
    input n1944;
    input n1943;
    input n1942;
    output ram_s_131_6;
    input n1941;
    output ram_s_131_5;
    input n1940;
    output ram_s_131_4;
    input n1939;
    output ram_s_131_3;
    input n1938;
    output ram_s_131_2;
    input n1937;
    output ram_s_131_1;
    input n1936;
    input n1935;
    input n1934;
    output ram_s_130_6;
    input n1933;
    output ram_s_130_5;
    input n1932;
    output ram_s_130_4;
    input n1931;
    output ram_s_130_3;
    input n1930;
    output ram_s_130_2;
    input n1929;
    output ram_s_130_1;
    input n1928;
    input n1927;
    input n1926;
    output ram_s_129_6;
    input n1925;
    output ram_s_129_5;
    input n1924;
    output ram_s_129_4;
    input n1923;
    output ram_s_129_3;
    input n1922;
    output ram_s_129_2;
    input n1921;
    output ram_s_129_1;
    input n1920;
    input n1919;
    input n1918;
    output ram_s_128_6;
    input n1917;
    output ram_s_128_5;
    input n1916;
    output ram_s_128_4;
    input n1915;
    output ram_s_128_3;
    input n1914;
    output ram_s_128_2;
    input n1913;
    output ram_s_128_1;
    input n1912;
    input n1543;
    output ram_s_81_7;
    input n1542;
    output ram_s_81_6;
    input n1541;
    input n1540;
    output ram_s_81_4;
    input n1539;
    output ram_s_81_3;
    input n1538;
    output ram_s_81_2;
    input n1537;
    output ram_s_81_1;
    input n1536;
    output ram_s_81_0;
    input n1495;
    input n1494;
    output ram_s_75_6;
    input n1493;
    output ram_s_75_5;
    input n1492;
    input n1491;
    output ram_s_75_3;
    input n1490;
    input n1489;
    output ram_s_75_1;
    input n1488;
    output ram_s_75_0;
    input n1487;
    input n1486;
    output ram_s_74_6;
    input n1485;
    output ram_s_74_5;
    input n1484;
    input n1483;
    output ram_s_74_3;
    input n1482;
    input n1481;
    output ram_s_74_1;
    input n1480;
    output ram_s_74_0;
    input n1479;
    input n1478;
    output ram_s_73_6;
    input n1477;
    output ram_s_73_5;
    input n1476;
    input n1475;
    output ram_s_73_3;
    input n1474;
    input n1473;
    output ram_s_73_1;
    input n1472;
    output ram_s_73_0;
    input n1471;
    input n1470;
    output ram_s_72_6;
    input n1469;
    output ram_s_72_5;
    input n1468;
    input n1467;
    output ram_s_72_3;
    input n1466;
    input n1465;
    output ram_s_72_1;
    input n1464;
    output ram_s_72_0;
    input n1463;
    output ram_s_71_7;
    input n1462;
    output ram_s_71_6;
    input n1461;
    output ram_s_71_5;
    input n1460;
    input n1459;
    input n1458;
    output ram_s_71_2;
    input n1457;
    output ram_s_71_1;
    input n1456;
    output ram_s_71_0;
    input n1455;
    output ram_s_70_7;
    input n1454;
    output ram_s_70_6;
    input n1453;
    output ram_s_70_5;
    input n1452;
    input n1451;
    input n1450;
    output ram_s_70_2;
    input n1449;
    output ram_s_70_1;
    input n1448;
    output ram_s_70_0;
    input n1447;
    output ram_s_69_7;
    input n1446;
    output ram_s_69_6;
    input n1445;
    output ram_s_69_5;
    input n1444;
    input n1443;
    input n1442;
    output ram_s_69_2;
    input n1441;
    output ram_s_69_1;
    input n1440;
    output ram_s_69_0;
    input n1439;
    output ram_s_68_7;
    input n1438;
    output ram_s_68_6;
    input n1437;
    output ram_s_68_5;
    input n1436;
    input n1435;
    input n1434;
    output ram_s_68_2;
    input n1433;
    output ram_s_68_1;
    input n1432;
    output ram_s_68_0;
    input n1431;
    output ram_s_67_7;
    input n1430;
    output ram_s_67_6;
    input n1429;
    output ram_s_67_5;
    input n1428;
    input n1427;
    output ram_s_67_3;
    input n1426;
    output ram_s_67_2;
    input n1425;
    output ram_s_67_1;
    input n1424;
    input n1423;
    output ram_s_66_7;
    input n1422;
    output ram_s_66_6;
    input n1421;
    output ram_s_66_5;
    input n1420;
    input n1419;
    output ram_s_66_3;
    input n1418;
    output ram_s_66_2;
    input n1417;
    output ram_s_66_1;
    input n1416;
    input n1415;
    output ram_s_65_7;
    input n1414;
    output ram_s_65_6;
    input n1413;
    output ram_s_65_5;
    input n1412;
    input n1411;
    output ram_s_65_3;
    input n1410;
    output ram_s_65_2;
    input n1409;
    output ram_s_65_1;
    input n1408;
    input n1407;
    output ram_s_64_7;
    input n1406;
    output ram_s_64_6;
    input n1405;
    output ram_s_64_5;
    input n1404;
    input n1403;
    output ram_s_64_3;
    input n1402;
    output ram_s_64_2;
    input n1401;
    output ram_s_64_1;
    input n1400;
    input n1399;
    output ram_s_63_7;
    input n1398;
    output ram_s_63_6;
    input n1397;
    output ram_s_63_5;
    input n1396;
    input n1395;
    output ram_s_63_3;
    input n1394;
    output ram_s_63_2;
    input n1393;
    output ram_s_63_1;
    input n1392;
    input n1391;
    output ram_s_62_7;
    input n1390;
    output ram_s_62_6;
    input n1389;
    output ram_s_62_5;
    input n1388;
    input n1387;
    output ram_s_62_3;
    input n1386;
    output ram_s_62_2;
    input n1385;
    output ram_s_62_1;
    input n1384;
    input n1359;
    output ram_s_58_7;
    input n1358;
    output ram_s_58_6;
    input n1357;
    input n1356;
    output ram_s_58_4;
    input n1355;
    output ram_s_58_3;
    input n1354;
    output ram_s_58_2;
    input n1353;
    output ram_s_58_1;
    input n1352;
    input n1351;
    output ram_s_57_7;
    input n1350;
    output ram_s_57_6;
    input n1349;
    input n1348;
    output ram_s_57_4;
    input n1347;
    output ram_s_57_3;
    input n1346;
    output ram_s_57_2;
    input n1345;
    output ram_s_57_1;
    input n1344;
    input n1271;
    output ram_s_47_7;
    input n1270;
    output ram_s_47_6;
    input n1269;
    output ram_s_47_5;
    input n1268;
    output ram_s_47_4;
    input n1267;
    output ram_s_47_3;
    input n1266;
    input n1265;
    output ram_s_47_1;
    input n1264;
    output ram_s_47_0;
    input n1255;
    output ram_s_45_7;
    input n1254;
    output ram_s_45_6;
    input n1253;
    output ram_s_45_5;
    input n1252;
    output ram_s_45_4;
    input n1251;
    output ram_s_45_3;
    input n1250;
    input n1249;
    output ram_s_45_1;
    input n1248;
    output ram_s_45_0;
    input n1247;
    output ram_s_44_7;
    input n1246;
    output ram_s_44_6;
    input n1245;
    output ram_s_44_5;
    input n1244;
    output ram_s_44_4;
    input n1243;
    output ram_s_44_3;
    input n1242;
    input n1241;
    output ram_s_44_1;
    input n1240;
    output ram_s_44_0;
    input n1239;
    input n1238;
    output ram_s_43_6;
    input n1237;
    output ram_s_43_5;
    input n1236;
    output ram_s_43_4;
    input n1235;
    output ram_s_43_3;
    input n1234;
    input n1233;
    input n1232;
    output ram_s_43_0;
    input n1215;
    input n1214;
    output ram_s_40_6;
    input n1213;
    output ram_s_40_5;
    input n1212;
    output ram_s_40_4;
    input n1211;
    output ram_s_40_3;
    input n1210;
    input n1209;
    input n1208;
    output ram_s_40_0;
    input n1207;
    input n1206;
    output ram_s_39_6;
    input n1205;
    output ram_s_39_5;
    input n1204;
    output ram_s_39_4;
    input n1203;
    output ram_s_39_3;
    input n1202;
    output ram_s_39_2;
    input n1201;
    output ram_s_39_1;
    input n1200;
    input n1199;
    input n1198;
    output ram_s_38_6;
    input n1197;
    output ram_s_38_5;
    input n1196;
    output ram_s_38_4;
    input n1195;
    output ram_s_38_3;
    input n1194;
    output ram_s_38_2;
    input n1193;
    output ram_s_38_1;
    input n1192;
    input n1191;
    input n1190;
    output ram_s_37_6;
    input n1189;
    output ram_s_37_5;
    input n1188;
    output ram_s_37_4;
    input n1187;
    output ram_s_37_3;
    input n1186;
    output ram_s_37_2;
    input n1185;
    output ram_s_37_1;
    input n1184;
    input n1183;
    input n1182;
    output ram_s_36_6;
    input n1181;
    output ram_s_36_5;
    input n1180;
    output ram_s_36_4;
    input n1179;
    output ram_s_36_3;
    input n1178;
    output ram_s_36_2;
    input n1177;
    output ram_s_36_1;
    input n1176;
    input n1175;
    input n1174;
    output ram_s_35_6;
    input n1173;
    output ram_s_35_5;
    input n1172;
    output ram_s_35_4;
    input n1171;
    output ram_s_35_3;
    input n1170;
    input n1169;
    input n1168;
    output ram_s_35_0;
    input n1167;
    input n1166;
    output ram_s_34_6;
    input n1165;
    output ram_s_34_5;
    input n1164;
    output ram_s_34_4;
    input n1163;
    output ram_s_34_3;
    input n1162;
    input n1161;
    input n1160;
    output ram_s_34_0;
    input n1159;
    input n1158;
    output ram_s_33_6;
    input n1157;
    output ram_s_33_5;
    input n1156;
    output ram_s_33_4;
    input n1155;
    output ram_s_33_3;
    input n1154;
    input n1153;
    input n1152;
    output ram_s_33_0;
    input n1151;
    input n1150;
    output ram_s_32_6;
    input n1149;
    output ram_s_32_5;
    input n1148;
    output ram_s_32_4;
    input n1147;
    output ram_s_32_3;
    input n1146;
    input n1145;
    input n1144;
    output ram_s_32_0;
    input n1051;
    input n1047;
    input n1046;
    input n1045;
    output ram_s_0_2;
    input n1044;
    output ram_s_12_3;
    input n1043;
    input n1042;
    output ram_s_11_1;
    input n1041;
    input n1040;
    output ram_s_12_1;
    input n1038;
    output ram_s_11_4;
    output n182;
    input n1037;
    output ram_s_12_4;
    output n54;
    input n1036;
    output ram_s_11_7;
    output n183;
    input n1035;
    output n55;
    input n1034;
    output ram_s_12_7;
    output n184;
    input n1033;
    output ram_s_12_2;
    output n56;
    input n1032;
    output ram_s_11_5;
    output n185;
    input n1031;
    output n57;
    input n1030;
    output ram_s_12_0;
    output n186;
    input n1029;
    output ram_s_11_3;
    output n58;
    output n187;
    output n59;
    output n188;
    output n60;
    output n189;
    output n61;
    output n190;
    output n62;
    output n191;
    output n63;
    output n192;
    input n1017;
    output ram_s_0_3;
    output n64;
    input n1016;
    output ram_s_0_4;
    output n193;
    input n1015;
    output ram_s_0_5;
    output n65;
    input n1014;
    output ram_s_0_6;
    output n194;
    input n1013;
    output n66;
    input n1012;
    output n195;
    input n1011;
    output n67;
    input n1010;
    output ram_s_1_2;
    input n1009;
    output ram_s_1_3;
    input n1008;
    output ram_s_1_4;
    input n1007;
    output ram_s_1_5;
    input n1006;
    output ram_s_4_4;
    input n1005;
    input n1004;
    input n1003;
    output ram_s_5_0;
    input n1002;
    output ram_s_4_6;
    input n1001;
    output ram_s_5_1;
    input n998;
    output ram_s_8_5;
    input n997;
    input n996;
    input n995;
    output ram_s_7_4;
    input n994;
    output ram_s_7_1;
    input n993;
    output ram_s_6_6;
    input n992;
    output ram_s_6_3;
    input n989;
    input n988;
    output ram_s_8_3;
    input n987;
    output ram_s_8_0;
    input n986;
    output n199;
    input n985;
    output ram_s_7_2;
    output n71;
    input n984;
    output n200;
    input n983;
    output ram_s_6_4;
    output n72;
    input n980;
    output ram_s_8_7;
    input n979;
    output ram_s_8_4;
    input n978;
    output ram_s_8_1;
    input n977;
    output ram_s_7_6;
    input n976;
    output ram_s_7_3;
    input n975;
    output ram_s_7_0;
    input n974;
    input n973;
    output ram_s_1_6;
    input n972;
    input n971;
    input n970;
    input n969;
    output ram_s_2_2;
    input n968;
    output ram_s_2_3;
    input n967;
    output ram_s_2_4;
    input n966;
    output ram_s_2_5;
    input n965;
    output ram_s_2_6;
    input n964;
    input n963;
    input n962;
    input n961;
    output ram_s_3_2;
    input n960;
    output ram_s_3_3;
    input n959;
    output ram_s_3_4;
    input n958;
    output ram_s_3_5;
    input n957;
    output ram_s_14_7;
    input n952;
    output ram_s_3_6;
    input n950;
    input n946;
    output ram_s_4_0;
    input n944;
    output ram_s_4_1;
    input n941;
    output ram_s_4_2;
    input n940;
    output ram_s_5_2;
    input n939;
    output ram_s_5_3;
    input n935;
    input n934;
    output ram_s_6_0;
    input n933;
    output ram_s_6_1;
    input n932;
    output ram_s_6_2;
    input n931;
    output ram_s_5_6;
    input n930;
    input n927;
    output ram_s_4_3;
    input n926;
    input n925;
    output ram_s_13_3;
    input n924;
    output ram_s_13_4;
    input n923;
    output n210;
    output n82;
    output n212;
    output n84;
    output n213;
    output n85;
    output n214;
    output n86;
    output n217;
    output n89;
    output n218;
    output n90;
    output n219;
    output n91;
    output n220;
    output n92;
    output n221;
    output n93;
    output n222;
    output n94;
    output n223;
    output n95;
    output n224;
    output n96;
    output n225;
    output n97;
    input n918;
    output ram_s_13_7;
    input n917;
    output ram_s_14_0;
    input n916;
    output ram_s_14_1;
    output n244;
    output n116;
    output n115;
    output n243;
    output n245;
    output n117;
    output n246;
    output n118;
    output n48;
    output n176;
    output n249;
    output n121;
    output n250;
    output n122;
    output n251;
    output n123;
    output n252;
    output n124;
    output n253;
    output n125;
    output n254;
    output n126;
    output n255;
    output n127;
    output n256;
    output n128;
    output n257;
    output n129;
    output ram_s_14_2;
    output ram_s_13_2;
    output ram_s_11_0;
    input n911;
    input n909;
    input n908;
    output ram_s_14_3;
    input n907;
    output ram_s_13_1;
    input n906;
    input n904;
    output ram_s_13_0;
    input n901;
    output ram_s_5_4;
    input n899;
    output LED1_c_0;
    input n765;
    input n938;
    output \pc_value[0] ;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [11:0]stack_memory;   // src/zipi8.vhd(322[13:25])
    wire [11:0]return_vector;   // src/x12_bit_program_address_generator.vhd(48[12:25])
    wire [11:0]pc_vector;   // src/zipi8.vhd(313[12:21])
    wire [7:0]alu_result;   // src/zipi8.vhd(344[12:22])
    wire [4:0]sx_addr;   // src/zipi8.vhd(286[12:19])
    wire [4:0]sy_addr;   // src/zipi8.vhd(287[12:19])
    
    wire register_enable;
    wire [11:0]register_vector;   // src/zipi8.vhd(312[12:27])
    
    wire t_state_2__N_28;
    wire [15:0]DI;   // src/ram.vhd(44[9:11])
    wire [4:0]stack_pointer_carry;   // src/zipi8.vhd(324[13:32])
    
    wire internal_reset_N_50, instruction_13_N_701, t_state_1_N_95, loadstar_type, 
        sx_addr4_value, shadow_zero_flag, shadow_bank, shadow_carry_flag, 
        pop_stack, push_stack_N_165, pop_stack_N_164;
    wire [11:0]address_c;   // src/top.vhd(80[20:27])
    wire [7:0]spm_data;   // src/zipi8.vhd(341[12:20])
    wire [7:0]port_id;   // src/zipi8.vhd(39[28:35])
    
    wire spm_enable;
    wire [7:0]shift_rotate_result;   // src/zipi8.vhd(338[12:31])
    
    wire flag_enable_type_N_217, regbank_type_N_77, n4283;
    wire [2:0]pc_mode;   // src/zipi8.vhd(293[12:19])
    wire [2:0]pc_mode_2__N_158;
    
    wire pc_mode_2__N_104, n6;
    wire [7:0]arith_logical_result;   // src/zipi8.vhd(334[12:32])
    wire [1:0]alu_mux_sel;   // src/zipi8.vhd(296[12:23])
    
    wire carry_arith_logical_7, carry_flag_value_N_436, flag_enable_type_N_216, 
        arith_carry_in;
    wire [1:0]alu_mux_sel_value;   // src/decode4alu.vhd(48[12:29])
    
    wire alu_mux_sel_value_0__N_184, arith_logical_sel_2__N_179, flag_enable;
    wire [2:0]arith_logical_sel;   // src/zipi8.vhd(297[12:29])
    
    wire n11080;
    wire [7:0]n409;
    
    wire n3783, n4, n11084;
    wire [7:0]half_arith_logical;   // src/arith_and_logic_operations.vhd(49[12:30])
    
    wire n722, n11107, n11109;
    wire [7:0]n417;
    
    wire n4_adj_885, n4247, flag_enable_type_N_222, pc_move_is_valid_o_N_132;
    
    x12_bit_program_address_generator x12_bit_program_address_generator_i (.stack_memory({stack_memory}), 
            .return_vector({Open_1, Open_2, Open_3, Open_4, Open_5, 
            Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, return_vector[0]}), 
            .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .\return_vector[3] (return_vector[3]), 
            .\return_vector[9] (return_vector[9]), .\instruction[1] (instruction[1]), 
            .\instruction[12] (instruction[12]), .\pc_vector[1] (pc_vector[1]), 
            .wea({wea}), .\instruction[2] (instruction[2]), .\pc_vector[2] (pc_vector[2]), 
            .\instruction[4] (instruction[4]), .\pc_vector[4] (pc_vector[4]), 
            .\instruction[5] (instruction[5]), .\pc_vector[5] (pc_vector[5]), 
            .\instruction[6] (instruction[6]), .\pc_vector[6] (pc_vector[6]), 
            .\instruction[11] (instruction[11]), .\pc_vector[11] (pc_vector[11]), 
            .\instruction[10] (instruction[10]), .\pc_vector[10] (pc_vector[10]), 
            .\instruction[8] (instruction[8]), .\pc_vector[8] (pc_vector[8]), 
            .\instruction[7] (instruction[7]), .\pc_vector[7] (pc_vector[7]));   // src/zipi8.vhd(446[42:75])
    two_banks_of_16_gp_reg two_banks_of_16_gp_reg_i (.CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), 
            .alu_result({alu_result}), .\sx_addr[4] (sx_addr[4]), .\instruction[11] (instruction[11]), 
            .\instruction[10] (instruction[10]), .\instruction[9] (instruction[9]), 
            .\instruction[8] (instruction[8]), .\sy_addr[4] (sy_addr[4]), 
            .\instruction[7] (instruction[7]), .\instruction[6] (instruction[6]), 
            .\instruction[5] (instruction[5]), .\instruction[4] (instruction[4]), 
            .register_enable(register_enable), .register_vector({\register_vector[11] , 
            \register_vector[10] , \register_vector[9] , \register_vector[8] , 
            register_vector[7:0]}), .\sx[7] (\sx[7] ), .\sx[6] (\sx[6] ), 
            .\sx[5] (\sx[5] ), .\sx[4] (\sx[4] ), .wea({wea}));   // src/zipi8.vhd(490[31:53])
    state_machine state_machine_i (.n8580(n8580), .bram_enable(bram_enable), 
            .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .\t_state[1] (\t_state[1] ), 
            .t_state_2__N_28(t_state_2__N_28), .internal_reset(internal_reset), 
            .BTN1_c(BTN1_c), .run(DI[3]), .\stack_pointer_carry[4] (stack_pointer_carry[4]), 
            .wea({wea}), .special_bit(special_bit), .internal_reset_N_50(internal_reset_N_50), 
            .\instruction[13] (instruction[13]), .instruction_13_N_701(instruction_13_N_701), 
            .t_state_1_N_95(t_state_1_N_95), .loadstar_type(loadstar_type), 
            .\sy_addr[4] (sy_addr[4]), .sx_addr4_value(sx_addr4_value));   // src/zipi8.vhd(354[22:35])
    stack stack_i (.CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .shadow_zero_flag(shadow_zero_flag), 
          .shadow_bank(shadow_bank), .special_bit(special_bit), .shadow_carry_flag(shadow_carry_flag), 
          .\stack_pointer_carry[4] (stack_pointer_carry[4]), .wea({wea}), 
          .bram_enable(bram_enable), .t_state_2__N_28(t_state_2__N_28), 
          .pop_stack(pop_stack), .\t_state[1] (\t_state[1] ), .internal_reset(internal_reset), 
          .t_state_1_N_95(t_state_1_N_95), .push_stack_N_165(push_stack_N_165), 
          .pop_stack_N_164(pop_stack_N_164), .\instruction[12] (instruction[12]), 
          .carry_flag(DI[0]), .zero_flag(DI[1]), .\sy_addr[4] (sy_addr[4]), 
          .run(DI[3]), .address({address_c[11], address[10:0]}), .VCC_net(VCC_net), 
          .stack_memory({stack_memory}));   // src/zipi8.vhd(470[14:19])
    spm_with_output_reg spm_with_output_reg_i (.spm_data({spm_data}), .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), 
            .port_id({port_id}), .ram_s_70_3(ram_s_70_3), .ram_s_71_3(ram_s_71_3), 
            .ram_s_69_3(ram_s_69_3), .ram_s_68_3(ram_s_68_3), .\sx[7] (\sx[7] ), 
            .\sx[6] (\sx[6] ), .\sx[5] (\sx[5] ), .\sx[4] (\sx[4] ), .\register_vector[10] (\register_vector[10] ), 
            .ram_s_34_7(ram_s_34_7), .ram_s_35_7(ram_s_35_7), .ram_s_33_7(ram_s_33_7), 
            .ram_s_32_7(ram_s_32_7), .\register_vector[9] (\register_vector[9] ), 
            .ram_s_11_6(ram_s_11_6), .ram_s_8_6(ram_s_8_6), .\register_vector[11] (\register_vector[11] ), 
            .ram_s_62_4(ram_s_62_4), .ram_s_63_4(ram_s_63_4), .ram_s_2_7(ram_s_2_7), 
            .ram_s_3_7(ram_s_3_7), .ram_s_1_7(ram_s_1_7), .ram_s_0_7(ram_s_0_7), 
            .ram_s_66_4(ram_s_66_4), .ram_s_67_4(ram_s_67_4), .ram_s_65_4(ram_s_65_4), 
            .ram_s_64_4(ram_s_64_4), .\register_vector[8] (\register_vector[8] ), 
            .ram_s_142_3(ram_s_142_3), .ram_s_141_3(ram_s_141_3), .ram_s_140_3(ram_s_140_3), 
            .ram_s_209_3(ram_s_209_3), .ram_s_130_0(ram_s_130_0), .ram_s_131_0(ram_s_131_0), 
            .ram_s_129_0(ram_s_129_0), .ram_s_128_0(ram_s_128_0), .ram_s_70_4(ram_s_70_4), 
            .ram_s_71_4(ram_s_71_4), .ram_s_69_4(ram_s_69_4), .ram_s_68_4(ram_s_68_4), 
            .ram_s_171_5(ram_s_171_5), .ram_s_168_5(ram_s_168_5), .ram_s_14_6(ram_s_14_6), 
            .ram_s_13_6(ram_s_13_6), .ram_s_12_6(ram_s_12_6), .ram_s_202_1(ram_s_202_1), 
            .ram_s_203_1(ram_s_203_1), .ram_s_6_5(ram_s_6_5), .ram_s_7_5(ram_s_7_5), 
            .ram_s_14_5(ram_s_14_5), .ram_s_5_5(ram_s_5_5), .ram_s_4_5(ram_s_4_5), 
            .ram_s_13_5(ram_s_13_5), .ram_s_12_5(ram_s_12_5), .ram_s_43_2(ram_s_43_2), 
            .ram_s_2_0(ram_s_2_0), .ram_s_3_0(ram_s_3_0), .ram_s_2_1(ram_s_2_1), 
            .ram_s_3_1(ram_s_3_1), .ram_s_1_0(ram_s_1_0), .ram_s_0_0(ram_s_0_0), 
            .ram_s_66_0(ram_s_66_0), .ram_s_67_0(ram_s_67_0), .ram_s_34_1(ram_s_34_1), 
            .ram_s_35_1(ram_s_35_1), .ram_s_33_1(ram_s_33_1), .ram_s_32_1(ram_s_32_1), 
            .ram_s_201_1(ram_s_201_1), .ram_s_200_1(ram_s_200_1), .ram_s_1_1(ram_s_1_1), 
            .ram_s_0_1(ram_s_0_1), .ram_s_65_0(ram_s_65_0), .ram_s_64_0(ram_s_64_0), 
            .ram_s_11_2(ram_s_11_2), .ram_s_8_2(ram_s_8_2), .ram_s_38_0(ram_s_38_0), 
            .ram_s_39_0(ram_s_39_0), .ram_s_40_2(ram_s_40_2), .ram_s_74_7(ram_s_74_7), 
            .ram_s_75_7(ram_s_75_7), .ram_s_73_7(ram_s_73_7), .ram_s_72_7(ram_s_72_7), 
            .ram_s_130_7(ram_s_130_7), .ram_s_131_7(ram_s_131_7), .ram_s_129_7(ram_s_129_7), 
            .ram_s_128_7(ram_s_128_7), .ram_s_37_0(ram_s_37_0), .ram_s_36_0(ram_s_36_0), 
            .ram_s_142_5(ram_s_142_5), .ram_s_141_5(ram_s_141_5), .ram_s_140_5(ram_s_140_5), 
            .ram_s_62_0(ram_s_62_0), .ram_s_63_0(ram_s_63_0), .ram_s_194_1(ram_s_194_1), 
            .ram_s_195_1(ram_s_195_1), .ram_s_193_1(ram_s_193_1), .ram_s_192_1(ram_s_192_1), 
            .ram_s_74_4(ram_s_74_4), .ram_s_75_4(ram_s_75_4), .ram_s_73_4(ram_s_73_4), 
            .ram_s_72_4(ram_s_72_4), .ram_s_43_7(ram_s_43_7), .ram_s_40_7(ram_s_40_7), 
            .ram_s_74_2(ram_s_74_2), .ram_s_75_2(ram_s_75_2), .ram_s_73_2(ram_s_73_2), 
            .ram_s_72_2(ram_s_72_2), .ram_s_186_3(ram_s_186_3), .ram_s_185_3(ram_s_185_3), 
            .ram_s_190_2(ram_s_190_2), .ram_s_191_2(ram_s_191_2), .ram_s_43_1(ram_s_43_1), 
            .wea({wea}), .ram_s_40_1(ram_s_40_1), .ram_s_6_7(ram_s_6_7), 
            .ram_s_7_7(ram_s_7_7), .ram_s_134_0(ram_s_134_0), .ram_s_135_0(ram_s_135_0), 
            .ram_s_5_7(ram_s_5_7), .ram_s_4_7(ram_s_4_7), .ram_s_133_0(ram_s_133_0), 
            .ram_s_132_0(ram_s_132_0), .ram_s_34_2(ram_s_34_2), .ram_s_35_2(ram_s_35_2), 
            .ram_s_58_5(ram_s_58_5), .ram_s_58_0(ram_s_58_0), .ram_s_57_0(ram_s_57_0), 
            .ram_s_139_0(ram_s_139_0), .ram_s_136_0(ram_s_136_0), .ram_s_190_5(ram_s_190_5), 
            .ram_s_191_5(ram_s_191_5), .ram_s_57_5(ram_s_57_5), .ram_s_33_2(ram_s_33_2), 
            .ram_s_32_2(ram_s_32_2), .ram_s_142_7(ram_s_142_7), .ram_s_141_7(ram_s_141_7), 
            .ram_s_140_7(ram_s_140_7), .ram_s_81_5(ram_s_81_5), .ram_s_190_1(ram_s_190_1), 
            .ram_s_191_1(ram_s_191_1), .ram_s_139_1(ram_s_139_1), .ram_s_136_1(ram_s_136_1), 
            .ram_s_38_7(ram_s_38_7), .ram_s_39_7(ram_s_39_7), .ram_s_37_7(ram_s_37_7), 
            .ram_s_36_7(ram_s_36_7), .n893(n893), .ram_s_14_4(ram_s_14_4), 
            .ram_s_190_7(ram_s_190_7), .ram_s_191_7(ram_s_191_7), .ram_s_47_2(ram_s_47_2), 
            .ram_s_45_2(ram_s_45_2), .ram_s_44_2(ram_s_44_2), .ram_s_134_5(ram_s_134_5), 
            .ram_s_135_5(ram_s_135_5), .ram_s_133_5(ram_s_133_5), .ram_s_132_5(ram_s_132_5), 
            .n2567(n2567), .ram_s_209_7(ram_s_209_7), .n2566(n2566), .ram_s_209_6(ram_s_209_6), 
            .n2565(n2565), .ram_s_209_5(ram_s_209_5), .n2564(n2564), .ram_s_209_4(ram_s_209_4), 
            .n2563(n2563), .n2562(n2562), .ram_s_209_2(ram_s_209_2), .n2561(n2561), 
            .ram_s_209_1(ram_s_209_1), .n2560(n2560), .ram_s_209_0(ram_s_209_0), 
            .n2519(n2519), .ram_s_203_7(ram_s_203_7), .n2518(n2518), .ram_s_203_6(ram_s_203_6), 
            .n2517(n2517), .ram_s_203_5(ram_s_203_5), .n2516(n2516), .ram_s_203_4(ram_s_203_4), 
            .n2515(n2515), .ram_s_203_3(ram_s_203_3), .n2514(n2514), .ram_s_203_2(ram_s_203_2), 
            .n2513(n2513), .n2512(n2512), .ram_s_203_0(ram_s_203_0), .n2511(n2511), 
            .ram_s_202_7(ram_s_202_7), .n2510(n2510), .ram_s_202_6(ram_s_202_6), 
            .n2509(n2509), .ram_s_202_5(ram_s_202_5), .n2508(n2508), .ram_s_202_4(ram_s_202_4), 
            .n2507(n2507), .ram_s_202_3(ram_s_202_3), .n2506(n2506), .ram_s_202_2(ram_s_202_2), 
            .n2505(n2505), .n2504(n2504), .ram_s_202_0(ram_s_202_0), .n2503(n2503), 
            .ram_s_201_7(ram_s_201_7), .n2502(n2502), .ram_s_201_6(ram_s_201_6), 
            .n2501(n2501), .ram_s_201_5(ram_s_201_5), .n2500(n2500), .ram_s_201_4(ram_s_201_4), 
            .n2499(n2499), .ram_s_201_3(ram_s_201_3), .n2498(n2498), .ram_s_201_2(ram_s_201_2), 
            .n2497(n2497), .n2496(n2496), .ram_s_201_0(ram_s_201_0), .n2495(n2495), 
            .ram_s_200_7(ram_s_200_7), .n2494(n2494), .ram_s_200_6(ram_s_200_6), 
            .n2493(n2493), .ram_s_200_5(ram_s_200_5), .n2492(n2492), .ram_s_200_4(ram_s_200_4), 
            .n2491(n2491), .ram_s_200_3(ram_s_200_3), .n2490(n2490), .ram_s_200_2(ram_s_200_2), 
            .n2489(n2489), .n2488(n2488), .ram_s_200_0(ram_s_200_0), .n2487(n2487), 
            .ram_s_199_7(ram_s_199_7), .n2486(n2486), .ram_s_199_6(ram_s_199_6), 
            .n2485(n2485), .ram_s_199_5(ram_s_199_5), .n2484(n2484), .ram_s_199_4(ram_s_199_4), 
            .n2483(n2483), .ram_s_199_3(ram_s_199_3), .n2482(n2482), .ram_s_199_2(ram_s_199_2), 
            .n2481(n2481), .ram_s_199_1(ram_s_199_1), .n2480(n2480), .ram_s_199_0(ram_s_199_0), 
            .n2479(n2479), .ram_s_198_7(ram_s_198_7), .n2478(n2478), .ram_s_198_6(ram_s_198_6), 
            .n2477(n2477), .ram_s_198_5(ram_s_198_5), .n2476(n2476), .ram_s_198_4(ram_s_198_4), 
            .n2475(n2475), .ram_s_198_3(ram_s_198_3), .n2474(n2474), .ram_s_198_2(ram_s_198_2), 
            .n2473(n2473), .ram_s_198_1(ram_s_198_1), .n2472(n2472), .ram_s_198_0(ram_s_198_0), 
            .n2471(n2471), .ram_s_197_7(ram_s_197_7), .n2470(n2470), .ram_s_197_6(ram_s_197_6), 
            .n2469(n2469), .ram_s_197_5(ram_s_197_5), .n2468(n2468), .ram_s_197_4(ram_s_197_4), 
            .n2467(n2467), .ram_s_197_3(ram_s_197_3), .n2466(n2466), .ram_s_197_2(ram_s_197_2), 
            .n2465(n2465), .ram_s_197_1(ram_s_197_1), .n2464(n2464), .ram_s_197_0(ram_s_197_0), 
            .n2463(n2463), .ram_s_196_7(ram_s_196_7), .n2462(n2462), .ram_s_196_6(ram_s_196_6), 
            .n2461(n2461), .ram_s_196_5(ram_s_196_5), .n2460(n2460), .ram_s_196_4(ram_s_196_4), 
            .n2459(n2459), .ram_s_196_3(ram_s_196_3), .n2458(n2458), .ram_s_196_2(ram_s_196_2), 
            .n2457(n2457), .ram_s_196_1(ram_s_196_1), .n2456(n2456), .ram_s_196_0(ram_s_196_0), 
            .n2455(n2455), .ram_s_195_7(ram_s_195_7), .n2454(n2454), .ram_s_195_6(ram_s_195_6), 
            .n2453(n2453), .ram_s_195_5(ram_s_195_5), .n2452(n2452), .ram_s_195_4(ram_s_195_4), 
            .n2451(n2451), .ram_s_195_3(ram_s_195_3), .n2450(n2450), .ram_s_195_2(ram_s_195_2), 
            .n2449(n2449), .n2448(n2448), .ram_s_195_0(ram_s_195_0), .n2447(n2447), 
            .ram_s_194_7(ram_s_194_7), .n2446(n2446), .ram_s_194_6(ram_s_194_6), 
            .n2445(n2445), .ram_s_194_5(ram_s_194_5), .n2444(n2444), .ram_s_194_4(ram_s_194_4), 
            .n2443(n2443), .ram_s_194_3(ram_s_194_3), .n2442(n2442), .ram_s_194_2(ram_s_194_2), 
            .n2441(n2441), .n2440(n2440), .ram_s_194_0(ram_s_194_0), .n2439(n2439), 
            .ram_s_193_7(ram_s_193_7), .n2438(n2438), .ram_s_193_6(ram_s_193_6), 
            .n2437(n2437), .ram_s_193_5(ram_s_193_5), .n2436(n2436), .ram_s_193_4(ram_s_193_4), 
            .n2435(n2435), .ram_s_193_3(ram_s_193_3), .n2434(n2434), .ram_s_193_2(ram_s_193_2), 
            .n2433(n2433), .n2432(n2432), .ram_s_193_0(ram_s_193_0), .n2431(n2431), 
            .ram_s_192_7(ram_s_192_7), .n2430(n2430), .ram_s_192_6(ram_s_192_6), 
            .n2429(n2429), .ram_s_192_5(ram_s_192_5), .n2428(n2428), .ram_s_192_4(ram_s_192_4), 
            .n2427(n2427), .ram_s_192_3(ram_s_192_3), .n2426(n2426), .ram_s_192_2(ram_s_192_2), 
            .n2425(n2425), .n2424(n2424), .ram_s_192_0(ram_s_192_0), .n2423(n2423), 
            .n2422(n2422), .ram_s_191_6(ram_s_191_6), .n2421(n2421), .n2420(n2420), 
            .ram_s_191_4(ram_s_191_4), .n2419(n2419), .ram_s_191_3(ram_s_191_3), 
            .n2418(n2418), .n2417(n2417), .n2416(n2416), .ram_s_191_0(ram_s_191_0), 
            .n2415(n2415), .n2414(n2414), .ram_s_190_6(ram_s_190_6), .n2413(n2413), 
            .n2412(n2412), .ram_s_190_4(ram_s_190_4), .n2411(n2411), .ram_s_190_3(ram_s_190_3), 
            .n2410(n2410), .n2409(n2409), .n2408(n2408), .ram_s_190_0(ram_s_190_0), 
            .n2383(n2383), .ram_s_186_7(ram_s_186_7), .n2382(n2382), .ram_s_186_6(ram_s_186_6), 
            .n2381(n2381), .ram_s_186_5(ram_s_186_5), .n2380(n2380), .ram_s_186_4(ram_s_186_4), 
            .n2379(n2379), .n2378(n2378), .ram_s_186_2(ram_s_186_2), .n2377(n2377), 
            .ram_s_186_1(ram_s_186_1), .n2376(n2376), .ram_s_186_0(ram_s_186_0), 
            .n2375(n2375), .ram_s_185_7(ram_s_185_7), .n2374(n2374), .ram_s_185_6(ram_s_185_6), 
            .n2373(n2373), .ram_s_185_5(ram_s_185_5), .n2372(n2372), .ram_s_185_4(ram_s_185_4), 
            .n2371(n2371), .n2370(n2370), .ram_s_185_2(ram_s_185_2), .n2369(n2369), 
            .ram_s_185_1(ram_s_185_1), .n2368(n2368), .ram_s_185_0(ram_s_185_0), 
            .n2295(n2295), .ram_s_175_7(ram_s_175_7), .n2294(n2294), .ram_s_175_6(ram_s_175_6), 
            .n2293(n2293), .ram_s_175_5(ram_s_175_5), .n2292(n2292), .ram_s_175_4(ram_s_175_4), 
            .n2291(n2291), .ram_s_175_3(ram_s_175_3), .n2290(n2290), .ram_s_175_2(ram_s_175_2), 
            .n2289(n2289), .ram_s_175_1(ram_s_175_1), .n2288(n2288), .ram_s_175_0(ram_s_175_0), 
            .n2279(n2279), .ram_s_173_7(ram_s_173_7), .n2278(n2278), .ram_s_173_6(ram_s_173_6), 
            .n2277(n2277), .ram_s_173_5(ram_s_173_5), .n2276(n2276), .ram_s_173_4(ram_s_173_4), 
            .n2275(n2275), .ram_s_173_3(ram_s_173_3), .n2274(n2274), .ram_s_173_2(ram_s_173_2), 
            .n2273(n2273), .ram_s_173_1(ram_s_173_1), .n2272(n2272), .ram_s_173_0(ram_s_173_0), 
            .n2271(n2271), .ram_s_172_7(ram_s_172_7), .n2270(n2270), .ram_s_172_6(ram_s_172_6), 
            .n2269(n2269), .ram_s_172_5(ram_s_172_5), .n2268(n2268), .ram_s_172_4(ram_s_172_4), 
            .n2267(n2267), .ram_s_172_3(ram_s_172_3), .n2266(n2266), .ram_s_172_2(ram_s_172_2), 
            .n2265(n2265), .ram_s_172_1(ram_s_172_1), .n2264(n2264), .ram_s_172_0(ram_s_172_0), 
            .n2263(n2263), .ram_s_171_7(ram_s_171_7), .n2262(n2262), .ram_s_171_6(ram_s_171_6), 
            .n2261(n2261), .n2260(n2260), .ram_s_171_4(ram_s_171_4), .n2259(n2259), 
            .ram_s_171_3(ram_s_171_3), .n2258(n2258), .ram_s_171_2(ram_s_171_2), 
            .n2257(n2257), .ram_s_171_1(ram_s_171_1), .n2256(n2256), .ram_s_171_0(ram_s_171_0), 
            .n2239(n2239), .ram_s_168_7(ram_s_168_7), .n2238(n2238), .ram_s_168_6(ram_s_168_6), 
            .n2237(n2237), .n2236(n2236), .ram_s_168_4(ram_s_168_4), .n2235(n2235), 
            .ram_s_168_3(ram_s_168_3), .n2234(n2234), .ram_s_168_2(ram_s_168_2), 
            .n2233(n2233), .ram_s_168_1(ram_s_168_1), .n2232(n2232), .ram_s_168_0(ram_s_168_0), 
            .n2231(n2231), .ram_s_167_7(ram_s_167_7), .n2230(n2230), .ram_s_167_6(ram_s_167_6), 
            .n2229(n2229), .ram_s_167_5(ram_s_167_5), .n2228(n2228), .ram_s_167_4(ram_s_167_4), 
            .n2227(n2227), .ram_s_167_3(ram_s_167_3), .n2226(n2226), .ram_s_167_2(ram_s_167_2), 
            .n2225(n2225), .ram_s_167_1(ram_s_167_1), .n2224(n2224), .ram_s_167_0(ram_s_167_0), 
            .n2223(n2223), .ram_s_166_7(ram_s_166_7), .n2222(n2222), .ram_s_166_6(ram_s_166_6), 
            .n2221(n2221), .ram_s_166_5(ram_s_166_5), .n2220(n2220), .ram_s_166_4(ram_s_166_4), 
            .n2219(n2219), .ram_s_166_3(ram_s_166_3), .n2218(n2218), .ram_s_166_2(ram_s_166_2), 
            .n2217(n2217), .ram_s_166_1(ram_s_166_1), .n2216(n2216), .ram_s_166_0(ram_s_166_0), 
            .n2215(n2215), .ram_s_165_7(ram_s_165_7), .n2214(n2214), .ram_s_165_6(ram_s_165_6), 
            .n2213(n2213), .ram_s_165_5(ram_s_165_5), .n2212(n2212), .ram_s_165_4(ram_s_165_4), 
            .n2211(n2211), .ram_s_165_3(ram_s_165_3), .n2210(n2210), .ram_s_165_2(ram_s_165_2), 
            .n2209(n2209), .ram_s_165_1(ram_s_165_1), .n2208(n2208), .ram_s_165_0(ram_s_165_0), 
            .n2207(n2207), .ram_s_164_7(ram_s_164_7), .n2206(n2206), .ram_s_164_6(ram_s_164_6), 
            .n2205(n2205), .ram_s_164_5(ram_s_164_5), .n2204(n2204), .ram_s_164_4(ram_s_164_4), 
            .n2203(n2203), .ram_s_164_3(ram_s_164_3), .n2202(n2202), .ram_s_164_2(ram_s_164_2), 
            .n2201(n2201), .ram_s_164_1(ram_s_164_1), .n2200(n2200), .ram_s_164_0(ram_s_164_0), 
            .n2199(n2199), .ram_s_163_7(ram_s_163_7), .n2198(n2198), .ram_s_163_6(ram_s_163_6), 
            .n2197(n2197), .ram_s_163_5(ram_s_163_5), .n2196(n2196), .ram_s_163_4(ram_s_163_4), 
            .n2195(n2195), .ram_s_163_3(ram_s_163_3), .n2194(n2194), .ram_s_163_2(ram_s_163_2), 
            .n2193(n2193), .ram_s_163_1(ram_s_163_1), .n2192(n2192), .ram_s_163_0(ram_s_163_0), 
            .n2191(n2191), .ram_s_162_7(ram_s_162_7), .n2190(n2190), .ram_s_162_6(ram_s_162_6), 
            .n2189(n2189), .ram_s_162_5(ram_s_162_5), .n2188(n2188), .ram_s_162_4(ram_s_162_4), 
            .n2187(n2187), .ram_s_162_3(ram_s_162_3), .n2186(n2186), .ram_s_162_2(ram_s_162_2), 
            .n2185(n2185), .ram_s_162_1(ram_s_162_1), .n2184(n2184), .ram_s_162_0(ram_s_162_0), 
            .n2183(n2183), .ram_s_161_7(ram_s_161_7), .n2182(n2182), .ram_s_161_6(ram_s_161_6), 
            .n2181(n2181), .ram_s_161_5(ram_s_161_5), .n2180(n2180), .ram_s_161_4(ram_s_161_4), 
            .n2179(n2179), .ram_s_161_3(ram_s_161_3), .n2178(n2178), .ram_s_161_2(ram_s_161_2), 
            .n2177(n2177), .ram_s_161_1(ram_s_161_1), .n2176(n2176), .ram_s_161_0(ram_s_161_0), 
            .n2175(n2175), .ram_s_160_7(ram_s_160_7), .n2174(n2174), .ram_s_160_6(ram_s_160_6), 
            .n2173(n2173), .ram_s_160_5(ram_s_160_5), .n2172(n2172), .ram_s_160_4(ram_s_160_4), 
            .n2171(n2171), .ram_s_160_3(ram_s_160_3), .n2170(n2170), .ram_s_160_2(ram_s_160_2), 
            .n2169(n2169), .ram_s_160_1(ram_s_160_1), .n2168(n2168), .ram_s_160_0(ram_s_160_0), 
            .n2031(n2031), .n2030(n2030), .ram_s_142_6(ram_s_142_6), .n2029(n2029), 
            .n2028(n2028), .ram_s_142_4(ram_s_142_4), .n2027(n2027), .n2026(n2026), 
            .ram_s_142_2(ram_s_142_2), .n2025(n2025), .ram_s_142_1(ram_s_142_1), 
            .n2024(n2024), .ram_s_142_0(ram_s_142_0), .n2023(n2023), .n2022(n2022), 
            .ram_s_141_6(ram_s_141_6), .n2021(n2021), .n2020(n2020), .ram_s_141_4(ram_s_141_4), 
            .n2019(n2019), .n2018(n2018), .ram_s_141_2(ram_s_141_2), .n2017(n2017), 
            .ram_s_141_1(ram_s_141_1), .n2016(n2016), .ram_s_141_0(ram_s_141_0), 
            .n2015(n2015), .n2014(n2014), .ram_s_140_6(ram_s_140_6), .n2013(n2013), 
            .n2012(n2012), .ram_s_140_4(ram_s_140_4), .n2011(n2011), .n2010(n2010), 
            .ram_s_140_2(ram_s_140_2), .n2009(n2009), .ram_s_140_1(ram_s_140_1), 
            .n2008(n2008), .ram_s_140_0(ram_s_140_0), .n2007(n2007), .ram_s_139_7(ram_s_139_7), 
            .n2006(n2006), .ram_s_139_6(ram_s_139_6), .n2005(n2005), .ram_s_139_5(ram_s_139_5), 
            .n2004(n2004), .ram_s_139_4(ram_s_139_4), .n2003(n2003), .ram_s_139_3(ram_s_139_3), 
            .n2002(n2002), .ram_s_139_2(ram_s_139_2), .n2001(n2001), .n2000(n2000), 
            .n1983(n1983), .ram_s_136_7(ram_s_136_7), .n1982(n1982), .ram_s_136_6(ram_s_136_6), 
            .n1981(n1981), .ram_s_136_5(ram_s_136_5), .n1980(n1980), .ram_s_136_4(ram_s_136_4), 
            .n1979(n1979), .ram_s_136_3(ram_s_136_3), .n1978(n1978), .ram_s_136_2(ram_s_136_2), 
            .n1977(n1977), .n1976(n1976), .n1975(n1975), .ram_s_135_7(ram_s_135_7), 
            .n1974(n1974), .ram_s_135_6(ram_s_135_6), .n1973(n1973), .n1972(n1972), 
            .ram_s_135_4(ram_s_135_4), .n1971(n1971), .ram_s_135_3(ram_s_135_3), 
            .n1970(n1970), .ram_s_135_2(ram_s_135_2), .n1969(n1969), .ram_s_135_1(ram_s_135_1), 
            .n1968(n1968), .n1967(n1967), .ram_s_134_7(ram_s_134_7), .n1966(n1966), 
            .ram_s_134_6(ram_s_134_6), .n1965(n1965), .n1964(n1964), .ram_s_134_4(ram_s_134_4), 
            .n1963(n1963), .ram_s_134_3(ram_s_134_3), .n1962(n1962), .ram_s_134_2(ram_s_134_2), 
            .n1961(n1961), .ram_s_134_1(ram_s_134_1), .n1960(n1960), .n1959(n1959), 
            .ram_s_133_7(ram_s_133_7), .n1958(n1958), .ram_s_133_6(ram_s_133_6), 
            .n1957(n1957), .n1956(n1956), .ram_s_133_4(ram_s_133_4), .n1955(n1955), 
            .ram_s_133_3(ram_s_133_3), .n1954(n1954), .ram_s_133_2(ram_s_133_2), 
            .n1953(n1953), .ram_s_133_1(ram_s_133_1), .n1952(n1952), .n1951(n1951), 
            .ram_s_132_7(ram_s_132_7), .n1950(n1950), .ram_s_132_6(ram_s_132_6), 
            .n1949(n1949), .n1948(n1948), .ram_s_132_4(ram_s_132_4), .n1947(n1947), 
            .ram_s_132_3(ram_s_132_3), .n1946(n1946), .ram_s_132_2(ram_s_132_2), 
            .n1945(n1945), .ram_s_132_1(ram_s_132_1), .n1944(n1944), .n1943(n1943), 
            .n1942(n1942), .ram_s_131_6(ram_s_131_6), .n1941(n1941), .ram_s_131_5(ram_s_131_5), 
            .n1940(n1940), .ram_s_131_4(ram_s_131_4), .n1939(n1939), .ram_s_131_3(ram_s_131_3), 
            .n1938(n1938), .ram_s_131_2(ram_s_131_2), .n1937(n1937), .ram_s_131_1(ram_s_131_1), 
            .n1936(n1936), .n1935(n1935), .n1934(n1934), .ram_s_130_6(ram_s_130_6), 
            .n1933(n1933), .ram_s_130_5(ram_s_130_5), .n1932(n1932), .ram_s_130_4(ram_s_130_4), 
            .n1931(n1931), .ram_s_130_3(ram_s_130_3), .n1930(n1930), .ram_s_130_2(ram_s_130_2), 
            .n1929(n1929), .ram_s_130_1(ram_s_130_1), .n1928(n1928), .n1927(n1927), 
            .n1926(n1926), .ram_s_129_6(ram_s_129_6), .n1925(n1925), .ram_s_129_5(ram_s_129_5), 
            .n1924(n1924), .ram_s_129_4(ram_s_129_4), .n1923(n1923), .ram_s_129_3(ram_s_129_3), 
            .n1922(n1922), .ram_s_129_2(ram_s_129_2), .n1921(n1921), .ram_s_129_1(ram_s_129_1), 
            .n1920(n1920), .n1919(n1919), .n1918(n1918), .ram_s_128_6(ram_s_128_6), 
            .n1917(n1917), .ram_s_128_5(ram_s_128_5), .n1916(n1916), .ram_s_128_4(ram_s_128_4), 
            .n1915(n1915), .ram_s_128_3(ram_s_128_3), .n1914(n1914), .ram_s_128_2(ram_s_128_2), 
            .n1913(n1913), .ram_s_128_1(ram_s_128_1), .n1912(n1912), .n1543(n1543), 
            .ram_s_81_7(ram_s_81_7), .n1542(n1542), .ram_s_81_6(ram_s_81_6), 
            .n1541(n1541), .n1540(n1540), .ram_s_81_4(ram_s_81_4), .n1539(n1539), 
            .ram_s_81_3(ram_s_81_3), .n1538(n1538), .ram_s_81_2(ram_s_81_2), 
            .n1537(n1537), .ram_s_81_1(ram_s_81_1), .n1536(n1536), .ram_s_81_0(ram_s_81_0), 
            .n1495(n1495), .n1494(n1494), .ram_s_75_6(ram_s_75_6), .n1493(n1493), 
            .ram_s_75_5(ram_s_75_5), .n1492(n1492), .n1491(n1491), .ram_s_75_3(ram_s_75_3), 
            .n1490(n1490), .n1489(n1489), .ram_s_75_1(ram_s_75_1), .n1488(n1488), 
            .ram_s_75_0(ram_s_75_0), .n1487(n1487), .n1486(n1486), .ram_s_74_6(ram_s_74_6), 
            .n1485(n1485), .ram_s_74_5(ram_s_74_5), .n1484(n1484), .n1483(n1483), 
            .ram_s_74_3(ram_s_74_3), .n1482(n1482), .n1481(n1481), .ram_s_74_1(ram_s_74_1), 
            .n1480(n1480), .ram_s_74_0(ram_s_74_0), .n1479(n1479), .n1478(n1478), 
            .ram_s_73_6(ram_s_73_6), .n1477(n1477), .ram_s_73_5(ram_s_73_5), 
            .n1476(n1476), .n1475(n1475), .ram_s_73_3(ram_s_73_3), .n1474(n1474), 
            .n1473(n1473), .ram_s_73_1(ram_s_73_1), .n1472(n1472), .ram_s_73_0(ram_s_73_0), 
            .n1471(n1471), .n1470(n1470), .ram_s_72_6(ram_s_72_6), .n1469(n1469), 
            .ram_s_72_5(ram_s_72_5), .n1468(n1468), .n1467(n1467), .ram_s_72_3(ram_s_72_3), 
            .n1466(n1466), .n1465(n1465), .ram_s_72_1(ram_s_72_1), .n1464(n1464), 
            .ram_s_72_0(ram_s_72_0), .n1463(n1463), .ram_s_71_7(ram_s_71_7), 
            .n1462(n1462), .ram_s_71_6(ram_s_71_6), .n1461(n1461), .ram_s_71_5(ram_s_71_5), 
            .n1460(n1460), .n1459(n1459), .n1458(n1458), .ram_s_71_2(ram_s_71_2), 
            .n1457(n1457), .ram_s_71_1(ram_s_71_1), .n1456(n1456), .ram_s_71_0(ram_s_71_0), 
            .n1455(n1455), .ram_s_70_7(ram_s_70_7), .n1454(n1454), .ram_s_70_6(ram_s_70_6), 
            .n1453(n1453), .ram_s_70_5(ram_s_70_5), .n1452(n1452), .n1451(n1451), 
            .n1450(n1450), .ram_s_70_2(ram_s_70_2), .n1449(n1449), .ram_s_70_1(ram_s_70_1), 
            .n1448(n1448), .ram_s_70_0(ram_s_70_0), .n1447(n1447), .ram_s_69_7(ram_s_69_7), 
            .n1446(n1446), .ram_s_69_6(ram_s_69_6), .n1445(n1445), .ram_s_69_5(ram_s_69_5), 
            .n1444(n1444), .n1443(n1443), .n1442(n1442), .ram_s_69_2(ram_s_69_2), 
            .n1441(n1441), .ram_s_69_1(ram_s_69_1), .n1440(n1440), .ram_s_69_0(ram_s_69_0), 
            .n1439(n1439), .ram_s_68_7(ram_s_68_7), .n1438(n1438), .ram_s_68_6(ram_s_68_6), 
            .n1437(n1437), .ram_s_68_5(ram_s_68_5), .n1436(n1436), .n1435(n1435), 
            .n1434(n1434), .ram_s_68_2(ram_s_68_2), .n1433(n1433), .ram_s_68_1(ram_s_68_1), 
            .n1432(n1432), .ram_s_68_0(ram_s_68_0), .n1431(n1431), .ram_s_67_7(ram_s_67_7), 
            .n1430(n1430), .ram_s_67_6(ram_s_67_6), .n1429(n1429), .ram_s_67_5(ram_s_67_5), 
            .n1428(n1428), .n1427(n1427), .ram_s_67_3(ram_s_67_3), .n1426(n1426), 
            .ram_s_67_2(ram_s_67_2), .n1425(n1425), .ram_s_67_1(ram_s_67_1), 
            .n1424(n1424), .n1423(n1423), .ram_s_66_7(ram_s_66_7), .n1422(n1422), 
            .ram_s_66_6(ram_s_66_6), .n1421(n1421), .ram_s_66_5(ram_s_66_5), 
            .n1420(n1420), .n1419(n1419), .ram_s_66_3(ram_s_66_3), .n1418(n1418), 
            .ram_s_66_2(ram_s_66_2), .n1417(n1417), .ram_s_66_1(ram_s_66_1), 
            .n1416(n1416), .n1415(n1415), .ram_s_65_7(ram_s_65_7), .n1414(n1414), 
            .ram_s_65_6(ram_s_65_6), .n1413(n1413), .ram_s_65_5(ram_s_65_5), 
            .n1412(n1412), .n1411(n1411), .ram_s_65_3(ram_s_65_3), .n1410(n1410), 
            .ram_s_65_2(ram_s_65_2), .n1409(n1409), .ram_s_65_1(ram_s_65_1), 
            .n1408(n1408), .n1407(n1407), .ram_s_64_7(ram_s_64_7), .n1406(n1406), 
            .ram_s_64_6(ram_s_64_6), .n1405(n1405), .ram_s_64_5(ram_s_64_5), 
            .n1404(n1404), .n1403(n1403), .ram_s_64_3(ram_s_64_3), .n1402(n1402), 
            .ram_s_64_2(ram_s_64_2), .n1401(n1401), .ram_s_64_1(ram_s_64_1), 
            .n1400(n1400), .n1399(n1399), .ram_s_63_7(ram_s_63_7), .n1398(n1398), 
            .ram_s_63_6(ram_s_63_6), .n1397(n1397), .ram_s_63_5(ram_s_63_5), 
            .n1396(n1396), .n1395(n1395), .ram_s_63_3(ram_s_63_3), .n1394(n1394), 
            .ram_s_63_2(ram_s_63_2), .n1393(n1393), .ram_s_63_1(ram_s_63_1), 
            .n1392(n1392), .n1391(n1391), .ram_s_62_7(ram_s_62_7), .n1390(n1390), 
            .ram_s_62_6(ram_s_62_6), .n1389(n1389), .ram_s_62_5(ram_s_62_5), 
            .n1388(n1388), .n1387(n1387), .ram_s_62_3(ram_s_62_3), .n1386(n1386), 
            .ram_s_62_2(ram_s_62_2), .n1385(n1385), .ram_s_62_1(ram_s_62_1), 
            .n1384(n1384), .n1359(n1359), .ram_s_58_7(ram_s_58_7), .n1358(n1358), 
            .ram_s_58_6(ram_s_58_6), .n1357(n1357), .n1356(n1356), .ram_s_58_4(ram_s_58_4), 
            .n1355(n1355), .ram_s_58_3(ram_s_58_3), .n1354(n1354), .ram_s_58_2(ram_s_58_2), 
            .n1353(n1353), .ram_s_58_1(ram_s_58_1), .n1352(n1352), .n1351(n1351), 
            .ram_s_57_7(ram_s_57_7), .n1350(n1350), .ram_s_57_6(ram_s_57_6), 
            .n1349(n1349), .n1348(n1348), .ram_s_57_4(ram_s_57_4), .n1347(n1347), 
            .ram_s_57_3(ram_s_57_3), .n1346(n1346), .ram_s_57_2(ram_s_57_2), 
            .n1345(n1345), .ram_s_57_1(ram_s_57_1), .n1344(n1344), .n1271(n1271), 
            .ram_s_47_7(ram_s_47_7), .n1270(n1270), .ram_s_47_6(ram_s_47_6), 
            .n1269(n1269), .ram_s_47_5(ram_s_47_5), .n1268(n1268), .ram_s_47_4(ram_s_47_4), 
            .n1267(n1267), .ram_s_47_3(ram_s_47_3), .n1266(n1266), .n1265(n1265), 
            .ram_s_47_1(ram_s_47_1), .n1264(n1264), .ram_s_47_0(ram_s_47_0), 
            .n1255(n1255), .ram_s_45_7(ram_s_45_7), .n1254(n1254), .ram_s_45_6(ram_s_45_6), 
            .n1253(n1253), .ram_s_45_5(ram_s_45_5), .n1252(n1252), .ram_s_45_4(ram_s_45_4), 
            .n1251(n1251), .ram_s_45_3(ram_s_45_3), .n1250(n1250), .n1249(n1249), 
            .ram_s_45_1(ram_s_45_1), .n1248(n1248), .ram_s_45_0(ram_s_45_0), 
            .n1247(n1247), .ram_s_44_7(ram_s_44_7), .n1246(n1246), .ram_s_44_6(ram_s_44_6), 
            .n1245(n1245), .ram_s_44_5(ram_s_44_5), .n1244(n1244), .ram_s_44_4(ram_s_44_4), 
            .n1243(n1243), .ram_s_44_3(ram_s_44_3), .n1242(n1242), .n1241(n1241), 
            .ram_s_44_1(ram_s_44_1), .n1240(n1240), .ram_s_44_0(ram_s_44_0), 
            .n1239(n1239), .n1238(n1238), .ram_s_43_6(ram_s_43_6), .n1237(n1237), 
            .ram_s_43_5(ram_s_43_5), .n1236(n1236), .ram_s_43_4(ram_s_43_4), 
            .n1235(n1235), .ram_s_43_3(ram_s_43_3), .n1234(n1234), .n1233(n1233), 
            .n1232(n1232), .ram_s_43_0(ram_s_43_0), .n1215(n1215), .n1214(n1214), 
            .ram_s_40_6(ram_s_40_6), .n1213(n1213), .ram_s_40_5(ram_s_40_5), 
            .n1212(n1212), .ram_s_40_4(ram_s_40_4), .n1211(n1211), .ram_s_40_3(ram_s_40_3), 
            .n1210(n1210), .n1209(n1209), .n1208(n1208), .ram_s_40_0(ram_s_40_0), 
            .n1207(n1207), .n1206(n1206), .ram_s_39_6(ram_s_39_6), .n1205(n1205), 
            .ram_s_39_5(ram_s_39_5), .n1204(n1204), .ram_s_39_4(ram_s_39_4), 
            .n1203(n1203), .ram_s_39_3(ram_s_39_3), .n1202(n1202), .ram_s_39_2(ram_s_39_2), 
            .n1201(n1201), .ram_s_39_1(ram_s_39_1), .n1200(n1200), .n1199(n1199), 
            .n1198(n1198), .ram_s_38_6(ram_s_38_6), .n1197(n1197), .ram_s_38_5(ram_s_38_5), 
            .n1196(n1196), .ram_s_38_4(ram_s_38_4), .n1195(n1195), .ram_s_38_3(ram_s_38_3), 
            .n1194(n1194), .ram_s_38_2(ram_s_38_2), .n1193(n1193), .ram_s_38_1(ram_s_38_1), 
            .n1192(n1192), .n1191(n1191), .n1190(n1190), .ram_s_37_6(ram_s_37_6), 
            .n1189(n1189), .ram_s_37_5(ram_s_37_5), .n1188(n1188), .ram_s_37_4(ram_s_37_4), 
            .n1187(n1187), .ram_s_37_3(ram_s_37_3), .n1186(n1186), .ram_s_37_2(ram_s_37_2), 
            .n1185(n1185), .ram_s_37_1(ram_s_37_1), .n1184(n1184), .n1183(n1183), 
            .n1182(n1182), .ram_s_36_6(ram_s_36_6), .n1181(n1181), .ram_s_36_5(ram_s_36_5), 
            .n1180(n1180), .ram_s_36_4(ram_s_36_4), .n1179(n1179), .ram_s_36_3(ram_s_36_3), 
            .n1178(n1178), .ram_s_36_2(ram_s_36_2), .n1177(n1177), .ram_s_36_1(ram_s_36_1), 
            .n1176(n1176), .n1175(n1175), .n1174(n1174), .ram_s_35_6(ram_s_35_6), 
            .n1173(n1173), .ram_s_35_5(ram_s_35_5), .n1172(n1172), .ram_s_35_4(ram_s_35_4), 
            .n1171(n1171), .ram_s_35_3(ram_s_35_3), .n1170(n1170), .n1169(n1169), 
            .n1168(n1168), .ram_s_35_0(ram_s_35_0), .n1167(n1167), .n1166(n1166), 
            .ram_s_34_6(ram_s_34_6), .n1165(n1165), .ram_s_34_5(ram_s_34_5), 
            .n1164(n1164), .ram_s_34_4(ram_s_34_4), .n1163(n1163), .ram_s_34_3(ram_s_34_3), 
            .n1162(n1162), .n1161(n1161), .n1160(n1160), .ram_s_34_0(ram_s_34_0), 
            .n1159(n1159), .n1158(n1158), .ram_s_33_6(ram_s_33_6), .n1157(n1157), 
            .ram_s_33_5(ram_s_33_5), .n1156(n1156), .ram_s_33_4(ram_s_33_4), 
            .n1155(n1155), .ram_s_33_3(ram_s_33_3), .n1154(n1154), .n1153(n1153), 
            .n1152(n1152), .ram_s_33_0(ram_s_33_0), .n1151(n1151), .n1150(n1150), 
            .ram_s_32_6(ram_s_32_6), .n1149(n1149), .ram_s_32_5(ram_s_32_5), 
            .n1148(n1148), .ram_s_32_4(ram_s_32_4), .n1147(n1147), .ram_s_32_3(ram_s_32_3), 
            .n1146(n1146), .n1145(n1145), .n1144(n1144), .ram_s_32_0(ram_s_32_0), 
            .n1051(n1051), .n1047(n1047), .n1046(n1046), .n1045(n1045), 
            .ram_s_0_2(ram_s_0_2), .n1044(n1044), .ram_s_12_3(ram_s_12_3), 
            .n1043(n1043), .n1042(n1042), .ram_s_11_1(ram_s_11_1), .n1041(n1041), 
            .n1040(n1040), .ram_s_12_1(ram_s_12_1), .n1038(n1038), .ram_s_11_4(ram_s_11_4), 
            .n182(n182), .n1037(n1037), .ram_s_12_4(ram_s_12_4), .n54(n54), 
            .n1036(n1036), .ram_s_11_7(ram_s_11_7), .n183(n183), .n1035(n1035), 
            .n55(n55), .n1034(n1034), .ram_s_12_7(ram_s_12_7), .n184(n184), 
            .n1033(n1033), .ram_s_12_2(ram_s_12_2), .n56(n56), .n1032(n1032), 
            .ram_s_11_5(ram_s_11_5), .n185(n185), .n1031(n1031), .n57(n57), 
            .n1030(n1030), .ram_s_12_0(ram_s_12_0), .n186(n186), .n1029(n1029), 
            .ram_s_11_3(ram_s_11_3), .n58(n58), .n187(n187), .n59(n59), 
            .n188(n188), .n60(n60), .n189(n189), .n61(n61), .n190(n190), 
            .n62(n62), .n191(n191), .n63(n63), .n192(n192), .n1017(n1017), 
            .ram_s_0_3(ram_s_0_3), .n64(n64), .n1016(n1016), .ram_s_0_4(ram_s_0_4), 
            .n193(n193), .n1015(n1015), .ram_s_0_5(ram_s_0_5), .n65(n65), 
            .n1014(n1014), .ram_s_0_6(ram_s_0_6), .n194(n194), .n1013(n1013), 
            .n66(n66), .n1012(n1012), .n195(n195), .n1011(n1011), .n67(n67), 
            .n1010(n1010), .ram_s_1_2(ram_s_1_2), .n1009(n1009), .ram_s_1_3(ram_s_1_3), 
            .n1008(n1008), .ram_s_1_4(ram_s_1_4), .n1007(n1007), .ram_s_1_5(ram_s_1_5), 
            .n1006(n1006), .ram_s_4_4(ram_s_4_4), .n1005(n1005), .n1004(n1004), 
            .n1003(n1003), .ram_s_5_0(ram_s_5_0), .n1002(n1002), .ram_s_4_6(ram_s_4_6), 
            .n1001(n1001), .ram_s_5_1(ram_s_5_1), .n998(n998), .ram_s_8_5(ram_s_8_5), 
            .n997(n997), .n996(n996), .n995(n995), .ram_s_7_4(ram_s_7_4), 
            .n994(n994), .ram_s_7_1(ram_s_7_1), .n993(n993), .ram_s_6_6(ram_s_6_6), 
            .n992(n992), .ram_s_6_3(ram_s_6_3), .n989(n989), .n988(n988), 
            .ram_s_8_3(ram_s_8_3), .n987(n987), .ram_s_8_0(ram_s_8_0), 
            .n986(n986), .n199(n199), .n985(n985), .ram_s_7_2(ram_s_7_2), 
            .n71(n71), .n984(n984), .n200(n200), .n983(n983), .ram_s_6_4(ram_s_6_4), 
            .n72(n72), .n980(n980), .ram_s_8_7(ram_s_8_7), .n979(n979), 
            .ram_s_8_4(ram_s_8_4), .n978(n978), .ram_s_8_1(ram_s_8_1), 
            .n977(n977), .ram_s_7_6(ram_s_7_6), .n976(n976), .ram_s_7_3(ram_s_7_3), 
            .n975(n975), .ram_s_7_0(ram_s_7_0), .n974(n974), .n973(n973), 
            .ram_s_1_6(ram_s_1_6), .n972(n972), .n971(n971), .n970(n970), 
            .n969(n969), .ram_s_2_2(ram_s_2_2), .n968(n968), .ram_s_2_3(ram_s_2_3), 
            .n967(n967), .ram_s_2_4(ram_s_2_4), .n966(n966), .ram_s_2_5(ram_s_2_5), 
            .n965(n965), .ram_s_2_6(ram_s_2_6), .n964(n964), .n963(n963), 
            .n962(n962), .n961(n961), .ram_s_3_2(ram_s_3_2), .n960(n960), 
            .ram_s_3_3(ram_s_3_3), .n959(n959), .ram_s_3_4(ram_s_3_4), 
            .n958(n958), .ram_s_3_5(ram_s_3_5), .n957(n957), .ram_s_14_7(ram_s_14_7), 
            .n952(n952), .ram_s_3_6(ram_s_3_6), .n950(n950), .n946(n946), 
            .ram_s_4_0(ram_s_4_0), .n944(n944), .ram_s_4_1(ram_s_4_1), 
            .n941(n941), .ram_s_4_2(ram_s_4_2), .n940(n940), .ram_s_5_2(ram_s_5_2), 
            .n939(n939), .ram_s_5_3(ram_s_5_3), .n935(n935), .n934(n934), 
            .ram_s_6_0(ram_s_6_0), .n933(n933), .ram_s_6_1(ram_s_6_1), 
            .n932(n932), .ram_s_6_2(ram_s_6_2), .n931(n931), .ram_s_5_6(ram_s_5_6), 
            .n930(n930), .n927(n927), .ram_s_4_3(ram_s_4_3), .n926(n926), 
            .n925(n925), .ram_s_13_3(ram_s_13_3), .n924(n924), .ram_s_13_4(ram_s_13_4), 
            .n923(n923), .n210(n210), .n82(n82), .n212(n212), .n84(n84), 
            .n213(n213), .n85(n85), .n214(n214), .n86(n86), .n217(n217), 
            .n89(n89), .n218(n218), .n90(n90), .n219(n219), .n91(n91), 
            .n220(n220), .n92(n92), .n221(n221), .n93(n93), .n222(n222), 
            .n94(n94), .n223(n223), .n95(n95), .n224(n224), .n96(n96), 
            .n225(n225), .n97(n97), .n918(n918), .ram_s_13_7(ram_s_13_7), 
            .n917(n917), .ram_s_14_0(ram_s_14_0), .n916(n916), .ram_s_14_1(ram_s_14_1), 
            .spm_enable(spm_enable), .n244(n244), .n116(n116), .n115(n115), 
            .n243(n243), .n245(n245), .n117(n117), .n246(n246), .n118(n118), 
            .n48(n48), .n176(n176), .n249(n249), .n121(n121), .n250(n250), 
            .n122(n122), .n251(n251), .n123(n123), .n252(n252), .n124(n124), 
            .n253(n253), .n125(n125), .n254(n254), .n126(n126), .n255(n255), 
            .n127(n127), .n256(n256), .n128(n128), .n257(n257), .n129(n129), 
            .ram_s_14_2(ram_s_14_2), .ram_s_13_2(ram_s_13_2), .ram_s_11_0(ram_s_11_0), 
            .n911(n911), .n909(n909), .n908(n908), .ram_s_14_3(ram_s_14_3), 
            .n907(n907), .ram_s_13_1(ram_s_13_1), .n906(n906), .n904(n904), 
            .ram_s_13_0(ram_s_13_0), .n901(n901), .ram_s_5_4(ram_s_5_4), 
            .n899(n899));   // src/zipi8.vhd(541[28:47])
    shift_and_rotate_operations shift_and_rotate_operations_i (.shift_rotate_result({shift_rotate_result}), 
            .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .\instruction[7] (instruction[7]), 
            .\sx[6] (\sx[6] ), .\instruction[3] (instruction[3]), .wea({wea}), 
            .\sx[5] (\sx[5] ), .\sx[7] (\sx[7] ), .\sx[4] (\sx[4] ), .\register_vector[11] (\register_vector[11] ), 
            .\register_vector[10] (\register_vector[10] ), .\register_vector[9] (\register_vector[9] ), 
            .\register_vector[8] (\register_vector[8] ), .\instruction[2] (instruction[2]), 
            .\instruction[0] (instruction[0]), .\instruction[1] (instruction[1]), 
            .carry_flag(DI[0]));   // src/zipi8.vhd(531[36:63])
    sel_of_out_port_value sel_of_out_port_value_i (.\register_vector[8] (\register_vector[8] ), 
            .\instruction[4] (instruction[4]), .\instruction[13] (instruction[13]), 
            .LED1_c_0(LED1_c_0), .wea({wea}));   // src/zipi8.vhd(512[30:51])
    sel_of_2nd_op_to_alu_and_port_id sel_of_2nd_op_to_alu_and_port_id_i (.\register_vector[7] (register_vector[7]), 
            .\instruction[7] (instruction[7]), .\instruction[12] (instruction[12]), 
            .port_id({port_id}), .wea({wea}), .\register_vector[2] (register_vector[2]), 
            .\instruction[2] (instruction[2]), .\register_vector[3] (register_vector[3]), 
            .\instruction[3] (instruction[3]), .\register_vector[4] (register_vector[4]), 
            .\instruction[4] (instruction[4]), .\register_vector[6] (register_vector[6]), 
            .\instruction[6] (instruction[6]), .\register_vector[5] (register_vector[5]), 
            .\instruction[5] (instruction[5]), .\register_vector[1] (register_vector[1]), 
            .\instruction[1] (instruction[1]), .\register_vector[0] (register_vector[0]), 
            .\instruction[0] (instruction[0]));   // src/zipi8.vhd(501[41:73])
    register_bank_control register_bank_control_i (.sx_addr4_value(sx_addr4_value), 
            .\sx_addr[4] (sx_addr[4]), .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .internal_reset_N_50(internal_reset_N_50), 
            .\sy_addr[4] (sy_addr[4]), .flag_enable_type_N_217(flag_enable_type_N_217), 
            .\instruction[16] (instruction[16]), .\instruction[14] (instruction[14]), 
            .\instruction[17] (instruction[17]), .loadstar_type(loadstar_type), 
            .regbank_type_N_77(regbank_type_N_77), .\instruction[15] (instruction[15]), 
            .n4283(n4283), .wea({wea}), .\instruction[12] (instruction[12]), 
            .\t_state[1] (\t_state[1] ), .shadow_bank(shadow_bank), .\instruction[0] (instruction[0]), 
            .internal_reset(internal_reset));   // src/zipi8.vhd(375[30:51])
    program_counter program_counter_i (.n765(n765), .address({address_c[11], 
            address[10:0]}), .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .internal_reset(internal_reset), 
            .n938(n938), .\pc_mode[0] (pc_mode[0]), .wea({wea}), .\pc_value[0] (\pc_value[0] ), 
            .\pc_vector[1] (pc_vector[1]), .register_vector({\register_vector[11] , 
            \register_vector[10] , \register_vector[9] , \register_vector[8] , 
            register_vector[7:0]}), .\instruction[0] (instruction[0]), .\return_vector[0] (return_vector[0]), 
            .\instruction[12] (instruction[12]), .\pc_vector[2] (pc_vector[2]), 
            .\pc_mode_2__N_158[2] (pc_mode_2__N_158[2]), .pc_mode_2__N_104(pc_mode_2__N_104), 
            .\instruction[3] (instruction[3]), .\return_vector[3] (return_vector[3]), 
            .\instruction[17] (instruction[17]), .\instruction[16] (instruction[16]), 
            .n6(n6), .\pc_vector[4] (pc_vector[4]), .\pc_vector[5] (pc_vector[5]), 
            .\pc_vector[6] (pc_vector[6]), .\pc_vector[11] (pc_vector[11]), 
            .\pc_vector[10] (pc_vector[10]), .\instruction[9] (instruction[9]), 
            .\return_vector[9] (return_vector[9]), .\pc_vector[8] (pc_vector[8]), 
            .\pc_vector[7] (pc_vector[7]));   // src/zipi8.vhd(457[24:39])
    mux_outputs_from_alu_spm_input_ports mux_outputs_from_alu_spm_input_ports_i (.arith_logical_result({arith_logical_result}), 
            .shift_rotate_result({shift_rotate_result}), .alu_mux_sel({alu_mux_sel}), 
            .wea({wea}), .spm_data({spm_data}), .alu_result({alu_result}));   // src/zipi8.vhd(550[46:82])
    flags flags_i (.CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .instruction_13_N_701(instruction_13_N_701), 
          .carry_arith_logical_7(carry_arith_logical_7), .zero_flag(DI[1]), 
          .internal_reset(internal_reset), .carry_flag(DI[0]), .\instruction[13] (instruction[13]), 
          .carry_flag_value_N_436(carry_flag_value_N_436), .flag_enable_type_N_216(flag_enable_type_N_216), 
          .arith_carry_in(arith_carry_in), .arith_logical_result({arith_logical_result}), 
          .wea({wea}), .\alu_mux_sel_value[1] (alu_mux_sel_value[1]), .alu_mux_sel_value_0__N_184(alu_mux_sel_value_0__N_184), 
          .\instruction[14] (instruction[14]), .arith_logical_sel_2__N_179(arith_logical_sel_2__N_179), 
          .flag_enable(flag_enable), .alu_result({alu_result}), .\instruction[15] (instruction[15]), 
          .\instruction[16] (instruction[16]), .shadow_zero_flag(shadow_zero_flag), 
          .\arith_logical_sel[0] (arith_logical_sel[0]), .\arith_logical_sel[2] (arith_logical_sel[2]), 
          .n11080(n11080), .\register_vector[9] (\register_vector[9] ), 
          .n338(n409[7]), .n3783(n3783), .n4(n4), .n11084(n11084), .\port_id[1] (port_id[1]), 
          .\half_arith_logical[1] (half_arith_logical[1]), .\sx[7] (\sx[7] ), 
          .\register_vector[8] (\register_vector[8] ), .\instruction[3] (instruction[3]), 
          .shadow_carry_flag(shadow_carry_flag), .\instruction[7] (instruction[7]), 
          .\port_id[5] (port_id[5]), .n722(n722), .n11107(n11107), .\sx[5] (\sx[5] ), 
          .n11109(n11109), .n350(n417[7]), .\half_arith_logical[5] (half_arith_logical[5]), 
          .n4_adj_2(n4_adj_885));   // src/zipi8.vhd(426[14:19])
    decode4alu decode4alu_i (.alu_mux_sel_value({alu_mux_sel_value[1], Open_12}), 
            .alu_mux_sel({alu_mux_sel}), .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), 
            .\instruction[16] (instruction[16]), .\instruction[15] (instruction[15]), 
            .\instruction[14] (instruction[14]), .carry_flag_value_N_436(carry_flag_value_N_436), 
            .wea({wea}), .alu_mux_sel_value_0__N_184(alu_mux_sel_value_0__N_184), 
            .arith_logical_sel({arith_logical_sel}), .n350(n417[7]), .n4247(n4247), 
            .arith_logical_sel_2__N_179(arith_logical_sel_2__N_179), .n722(n722), 
            .\instruction[13] (instruction[13]), .\sx[5] (\sx[5] ), .n338(n409[7]), 
            .n11109(n11109));   // src/zipi8.vhd(400[19:29])
    decode4_strobes_enables decode4_strobes_enables_i (.flag_enable(flag_enable), 
            .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .t_state_1_N_95(t_state_1_N_95), 
            .register_enable(register_enable), .spm_enable(spm_enable), 
            .instruction_13_N_701(instruction_13_N_701), .\instruction[17] (instruction[17]), 
            .\instruction[15] (instruction[15]), .\instruction[14] (instruction[14]), 
            .flag_enable_type_N_222(flag_enable_type_N_222), .wea({wea}), 
            .carry_flag(DI[0]), .pc_move_is_valid_o_N_132(pc_move_is_valid_o_N_132), 
            .\t_state[1] (\t_state[1] ), .arith_logical_sel_2__N_179(arith_logical_sel_2__N_179), 
            .\instruction[16] (instruction[16]), .flag_enable_type_N_216(flag_enable_type_N_216), 
            .n4247(n4247), .n4283(n4283), .\instruction[12] (instruction[12]), 
            .\instruction[13] (instruction[13]), .flag_enable_type_N_217(flag_enable_type_N_217));   // src/zipi8.vhd(410[32:55])
    decode4_pc_statck decode4_pc_statck_i (.\instruction[15] (instruction[15]), 
            .pc_mode_2__N_104(pc_mode_2__N_104), .\instruction[14] (instruction[14]), 
            .\instruction[12] (instruction[12]), .n6(n6), .regbank_type_N_77(regbank_type_N_77), 
            .\pc_mode_2__N_158[2] (pc_mode_2__N_158[2]), .pop_stack_N_164(pop_stack_N_164), 
            .push_stack_N_165(push_stack_N_165), .wea({wea}), .pop_stack(pop_stack), 
            .\instruction[17] (instruction[17]), .zero_flag(DI[1]), .pc_move_is_valid_o_N_132(pc_move_is_valid_o_N_132), 
            .flag_enable_type_N_222(flag_enable_type_N_222), .carry_flag(DI[0]), 
            .\instruction[13] (instruction[13]), .\instruction[16] (instruction[16]), 
            .n4283(n4283), .\pc_mode[0] (pc_mode[0]), .arith_logical_sel_2__N_179(arith_logical_sel_2__N_179));   // src/zipi8.vhd(389[26:43])
    arith_and_logic_operations arith_and_logic_operations_i (.arith_logical_result({arith_logical_result}), 
            .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .arith_logical_sel({arith_logical_sel}), 
            .\register_vector[8] (\register_vector[8] ), .n722(n722), .n4(n4), 
            .n11080(n11080), .arith_carry_in(arith_carry_in), .wea({wea}), 
            .\port_id[0] (port_id[0]), .\register_vector[10] (\register_vector[10] ), 
            .\port_id[2] (port_id[2]), .\half_arith_logical[1] (half_arith_logical[1]), 
            .\register_vector[9] (\register_vector[9] ), .\register_vector[11] (\register_vector[11] ), 
            .\port_id[3] (port_id[3]), .\sx[4] (\sx[4] ), .\port_id[4] (port_id[4]), 
            .\sx[6] (\sx[6] ), .\port_id[6] (port_id[6]), .\half_arith_logical[5] (half_arith_logical[5]), 
            .\sx[5] (\sx[5] ), .\sx[7] (\sx[7] ), .carry_arith_logical_7(carry_arith_logical_7), 
            .n350(n417[7]), .\port_id[7] (port_id[7]), .n11084(n11084), 
            .n3783(n3783), .\port_id[1] (port_id[1]), .n4247(n4247), .\instruction[14] (instruction[14]), 
            .n338(n409[7]), .n4_adj_1(n4_adj_885), .n11107(n11107));   // src/zipi8.vhd(520[36:62])
    
endmodule
//
// Verilog Description of module x12_bit_program_address_generator
//

module x12_bit_program_address_generator (stack_memory, return_vector, CLK_3P3_MHZ_c, 
            \return_vector[3] , \return_vector[9] , \instruction[1] , 
            \instruction[12] , \pc_vector[1] , wea, \instruction[2] , 
            \pc_vector[2] , \instruction[4] , \pc_vector[4] , \instruction[5] , 
            \pc_vector[5] , \instruction[6] , \pc_vector[6] , \instruction[11] , 
            \pc_vector[11] , \instruction[10] , \pc_vector[10] , \instruction[8] , 
            \pc_vector[8] , \instruction[7] , \pc_vector[7] );
    input [11:0]stack_memory;
    output [11:0]return_vector;
    input CLK_3P3_MHZ_c;
    output \return_vector[3] ;
    output \return_vector[9] ;
    input \instruction[1] ;
    input \instruction[12] ;
    output \pc_vector[1] ;
    input [0:0]wea;
    input \instruction[2] ;
    output \pc_vector[2] ;
    input \instruction[4] ;
    output \pc_vector[4] ;
    input \instruction[5] ;
    output \pc_vector[5] ;
    input \instruction[6] ;
    output \pc_vector[6] ;
    input \instruction[11] ;
    output \pc_vector[11] ;
    input \instruction[10] ;
    output \pc_vector[10] ;
    input \instruction[8] ;
    output \pc_vector[8] ;
    input \instruction[7] ;
    output \pc_vector[7] ;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [11:0]return_vector_c;   // src/x12_bit_program_address_generator.vhd(48[12:25])
    
    SB_DFF return_vector_i0 (.Q(return_vector[0]), .C(CLK_3P3_MHZ_c), .D(stack_memory[0]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i1 (.Q(return_vector_c[1]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[1]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i2 (.Q(return_vector_c[2]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[2]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i3 (.Q(\return_vector[3] ), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[3]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i4 (.Q(return_vector_c[4]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[4]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i5 (.Q(return_vector_c[5]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[5]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i6 (.Q(return_vector_c[6]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[6]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i7 (.Q(return_vector_c[7]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[7]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i8 (.Q(return_vector_c[8]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[8]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i9 (.Q(\return_vector[9] ), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[9]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i10 (.Q(return_vector_c[10]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[10]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_DFF return_vector_i11 (.Q(return_vector_c[11]), .C(CLK_3P3_MHZ_c), 
           .D(stack_memory[11]));   // src/x12_bit_program_address_generator.vhd(54[9] 56[16])
    SB_LUT4 i12_3_lut (.I0(\instruction[1] ), .I1(return_vector_c[1]), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(\pc_vector[1] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_3_lut (.I0(\instruction[2] ), .I1(return_vector_c[2]), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(\pc_vector[2] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15_3_lut (.I0(\instruction[4] ), .I1(return_vector_c[4]), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(\pc_vector[4] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_3_lut (.I0(\instruction[5] ), .I1(return_vector_c[5]), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(\pc_vector[5] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17_3_lut (.I0(\instruction[6] ), .I1(return_vector_c[6]), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(\pc_vector[6] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut (.I0(\instruction[11] ), .I1(return_vector_c[11]), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(\pc_vector[11] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21_3_lut (.I0(\instruction[10] ), .I1(return_vector_c[10]), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(\pc_vector[10] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_3_lut (.I0(\instruction[8] ), .I1(return_vector_c[8]), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(\pc_vector[8] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_3_lut (.I0(\instruction[7] ), .I1(return_vector_c[7]), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(\pc_vector[7] ));   // src/x12_bit_program_address_generator.vhd(235[25] 236[76])
    defparam i18_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module two_banks_of_16_gp_reg
//

module two_banks_of_16_gp_reg (CLK_3P3_MHZ_c, alu_result, \sx_addr[4] , 
            \instruction[11] , \instruction[10] , \instruction[9] , \instruction[8] , 
            \sy_addr[4] , \instruction[7] , \instruction[6] , \instruction[5] , 
            \instruction[4] , register_enable, register_vector, \sx[7] , 
            \sx[6] , \sx[5] , \sx[4] , wea);
    input CLK_3P3_MHZ_c;
    input [7:0]alu_result;
    input \sx_addr[4] ;
    input \instruction[11] ;
    input \instruction[10] ;
    input \instruction[9] ;
    input \instruction[8] ;
    input \sy_addr[4] ;
    input \instruction[7] ;
    input \instruction[6] ;
    input \instruction[5] ;
    input \instruction[4] ;
    input register_enable;
    output [11:0]register_vector;
    output \sx[7] ;
    output \sx[6] ;
    output \sx[5] ;
    output \sx[4] ;
    input [0:0]wea;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    ram32m_behav sy_bank (.WCLK(CLK_3P3_MHZ_c), .WE(register_enable), .DI({alu_result}), 
            .ADDR_RD({\sy_addr[4] , \instruction[7] , \instruction[6] , 
            \instruction[5] , \instruction[4] }), .ADDR_WR({\sx_addr[4] , 
            \instruction[11] , \instruction[10] , \instruction[9] , \instruction[8] }), 
            .DO({register_vector[7:0]})) /* synthesis LSE_LINE_FILE_ID=76, LSE_LCOL=31, LSE_RCOL=53, LSE_LLINE=490, LSE_RLINE=490 */ ;   // src/two_banks_of_16_gp_reg.vhd(151[14:26])
    defparam sy_bank.DATA_WIDTH = 8;
    defparam sy_bank.ADDRESS_WIDTH = 5;
    \ram(8,5)  sx_bank (.\instruction[9] (\instruction[9] ), .\instruction[10] (\instruction[10] ), 
            .\instruction[8] (\instruction[8] ), .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), 
            .\instruction[11] (\instruction[11] ), .\sx[7] (\sx[7] ), .\sx[6] (\sx[6] ), 
            .\sx[5] (\sx[5] ), .\sx[4] (\sx[4] ), .\register_vector[11] (register_vector[11]), 
            .\register_vector[10] (register_vector[10]), .\register_vector[9] (register_vector[9]), 
            .\register_vector[8] (register_vector[8]), .\sx_addr[4] (\sx_addr[4] ), 
            .alu_result({alu_result}), .wea({wea}), .register_enable(register_enable));   // src/two_banks_of_16_gp_reg.vhd(138[14:17])
    
endmodule
//
// Verilog Description of module ram32m_behav
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \ram(8,5) 
//

module \ram(8,5)  (\instruction[9] , \instruction[10] , \instruction[8] , 
            CLK_3P3_MHZ_c, \instruction[11] , \sx[7] , \sx[6] , \sx[5] , 
            \sx[4] , \register_vector[11] , \register_vector[10] , \register_vector[9] , 
            \register_vector[8] , \sx_addr[4] , alu_result, wea, register_enable);
    input \instruction[9] ;
    input \instruction[10] ;
    input \instruction[8] ;
    input CLK_3P3_MHZ_c;
    input \instruction[11] ;
    output \sx[7] ;
    output \sx[6] ;
    output \sx[5] ;
    output \sx[4] ;
    output \register_vector[11] ;
    output \register_vector[10] ;
    output \register_vector[9] ;
    output \register_vector[8] ;
    input \sx_addr[4] ;
    input [7:0]alu_result;
    input [0:0]wea;
    input register_enable;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    wire n11037, n11038, n11231, n11026, n11025, n11234, ram_s_26_6, 
        ram_s_27_6, n12365, ram_s_2_4, ram_s_3_4, n11519, ram_s_25_6, 
        ram_s_24_6, n12368, ram_s_1_4, ram_s_0_4, n11522, ram_s_10_2, 
        ram_s_11_2, n13037, ram_s_30_3, ram_s_31_3, n12131, ram_s_9_2, 
        ram_s_8_2, n13040, ram_s_29_3, ram_s_28_3, n12134, ram_s_30_0, 
        ram_s_31_0, n11927, ram_s_29_0, ram_s_28_0, n11012, n3192, 
        ram_s_31_7, n3191, ram_s_31_6, ram_s_18_0, ram_s_19_0, n11741, 
        ram_s_17_0, ram_s_16_0, n11744, n3190, ram_s_31_5, n3189, 
        ram_s_31_4, n3188, n3187, ram_s_31_2, n3186, ram_s_31_1, 
        n3185, n11846, n11828, n11915, n11882, n11900, n11918, 
        ram_s_26_2, ram_s_27_2, n12101, ram_s_30_7, n12995, n3184, 
        n3183, ram_s_30_6, n3182, ram_s_30_5, n3181, ram_s_30_4, 
        ram_s_29_7, ram_s_28_7, n10421, ram_s_25_2, ram_s_24_2, n8858, 
        n3180, ram_s_14_2, ram_s_15_2, n12977, ram_s_13_2, ram_s_12_2, 
        n12980, n3179, ram_s_30_2, n3178, ram_s_30_1, n3177, n3176, 
        n3174, ram_s_29_6, n3173, ram_s_29_5, n3172, ram_s_29_4, 
        n3171, n3170, ram_s_29_2, n3169, ram_s_29_1, n3168, n11492, 
        n11903, n3167, n11498, n11906, n3166, ram_s_28_6, n3165, 
        ram_s_28_5, n3164, ram_s_28_4, n3163, n3162, ram_s_28_2, 
        n3161, ram_s_28_1, n3160, n3159, ram_s_27_7, n3158, n3157, 
        ram_s_27_5, n3156, ram_s_27_4, n3155, ram_s_27_3, n3154, 
        n3153, ram_s_27_1, n3152, ram_s_27_0, n3151, ram_s_26_7, 
        n3150, n3149, ram_s_26_5, n3148, ram_s_26_4, n3147, ram_s_26_3, 
        n3146, n3145, ram_s_26_1, n3144, ram_s_26_0, n3143, ram_s_25_7, 
        n3142, n3141, ram_s_25_5, n3140, ram_s_25_4, n3139, ram_s_25_3, 
        n3138, n3137, ram_s_25_1, n3136, ram_s_25_0, n3135, ram_s_24_7, 
        n3134, n3133, ram_s_24_5, n3132, ram_s_24_4, n3131, ram_s_24_3, 
        n3130, n3129, ram_s_24_1, n3128, ram_s_24_0, n3127, ram_s_23_7, 
        n3126, ram_s_23_6, n3125, ram_s_23_5, ram_s_22_0, ram_s_23_0, 
        n11495, ram_s_2_0, ram_s_3_0, n11897, ram_s_21_0, ram_s_20_0, 
        n3124, ram_s_23_4, n3123, ram_s_23_3, n3122, ram_s_23_2, 
        n3121, ram_s_23_1, n3120, n3119, ram_s_22_7, n3118, ram_s_22_6, 
        n3117, ram_s_22_5, n3116, ram_s_22_4, ram_s_1_0, ram_s_0_0, 
        n11489, n3115, ram_s_22_3, n3114, ram_s_22_2, n3113, ram_s_22_1, 
        n3112, n3111, ram_s_21_7, n3110, ram_s_21_6, n3109, ram_s_21_5, 
        n3108, ram_s_21_4, ram_s_18_2, ram_s_19_2, n12923, n3107, 
        ram_s_21_3, n3106, ram_s_21_2, n3105, ram_s_21_1, n3104, 
        n3103, ram_s_20_7, n3102, ram_s_20_6, n3101, ram_s_20_5, 
        n3100, ram_s_20_4, n3099, ram_s_20_3, n3098, ram_s_20_2, 
        n3097, ram_s_20_1, n3096, n3095, ram_s_19_7, n3094, ram_s_19_6, 
        n3093, ram_s_19_5, n3092, ram_s_19_4, n3091, ram_s_19_3, 
        n3090, n3089, ram_s_19_1, n3088, n3087, ram_s_18_7, n3086, 
        ram_s_18_6, n3085, ram_s_18_5, ram_s_17_2, ram_s_16_2, n8840, 
        n3084, ram_s_18_4, n3083, ram_s_18_3, n3082, n3081, ram_s_18_1, 
        n3080, n3079, ram_s_17_7, n3078, ram_s_17_6, n3077, ram_s_17_5, 
        n3076, ram_s_17_4, n3075, ram_s_17_3, n3074, n3073, ram_s_17_1, 
        n3072, n3071, ram_s_16_7, n3070, ram_s_16_6, n3069, ram_s_16_5, 
        n3068, ram_s_16_4, n3067, ram_s_16_3, n3066, n3065, ram_s_16_1, 
        n3064, n3063, ram_s_15_7, n3062, ram_s_15_6, n3061, ram_s_15_5, 
        n3060, ram_s_15_4, n3059, ram_s_15_3, n3058, n3057, ram_s_15_1, 
        n3056, ram_s_15_0, n3055, ram_s_14_7, n3054, ram_s_14_6, 
        n3053, ram_s_14_5, n3052, ram_s_14_4, n3051, ram_s_14_3, 
        n3050, n3049, ram_s_14_1, n3048, ram_s_14_0, n3047, ram_s_13_7, 
        n3046, ram_s_13_6, n3045, ram_s_13_5, n3044, ram_s_13_4, 
        n3043, ram_s_13_3, n3042, n3041, ram_s_13_1, n3040, ram_s_13_0, 
        n3039, ram_s_12_7, n3038, ram_s_12_6, n3037, ram_s_12_5, 
        n3036, ram_s_12_4, n3035, ram_s_12_3, n3034, n3033, ram_s_12_1, 
        n3032, ram_s_12_0, n3031, ram_s_11_7, n3030, ram_s_11_6, 
        n3029, ram_s_11_5, n3028, ram_s_11_4, n3027, ram_s_11_3, 
        n3026, n3025, ram_s_11_1, n3024, ram_s_11_0, n3023, ram_s_10_7, 
        n3022, ram_s_10_6, n3021, ram_s_10_5, n3020, ram_s_10_4, 
        n3019, ram_s_10_3, n3018, n3017, ram_s_10_1, n3016, ram_s_10_0, 
        n3015, ram_s_9_7, n3014, ram_s_9_6, n3013, ram_s_9_5, n3012, 
        ram_s_9_4, n3011, ram_s_9_3, n3010, n3009, ram_s_9_1, n3008, 
        ram_s_9_0, n3007, ram_s_8_7, n3006, ram_s_8_6, n3005, ram_s_8_5, 
        n3004, ram_s_8_4, n3003, ram_s_8_3, n3002, n3001, ram_s_8_1, 
        n3000, ram_s_8_0, n2999, ram_s_7_7, n2998, ram_s_7_6, n2997, 
        ram_s_7_5, n2996, ram_s_7_4, n2995, ram_s_7_3, n2994, ram_s_7_2, 
        n2993, ram_s_7_1, n2992, ram_s_7_0, n2991, ram_s_6_7, n2990, 
        ram_s_6_6, n2989, ram_s_6_5, n2988, ram_s_6_4, n2987, ram_s_6_3, 
        n2986, ram_s_6_2, n2985, ram_s_6_1, n2984, ram_s_6_0, n2983, 
        ram_s_5_7, n2982, ram_s_5_6, n2981, ram_s_5_5, n2980, ram_s_5_4, 
        n2979, ram_s_5_3, n2978, ram_s_5_2, n2977, ram_s_5_1, n2976, 
        ram_s_5_0, n2975, ram_s_4_7, n2974, ram_s_4_6, n2973, ram_s_4_5, 
        n2972, ram_s_4_4, n2971, ram_s_4_3, n2970, ram_s_4_2, n2969, 
        ram_s_4_1, n2968, ram_s_4_0, n2967, ram_s_3_7, n2966, ram_s_3_6, 
        n2965, ram_s_3_5, n2964, n2963, ram_s_3_3, n2962, ram_s_3_2, 
        n2961, ram_s_3_1, n2960, n2959, ram_s_2_7, n2958, ram_s_2_6, 
        n2957, ram_s_2_5, n2956, n2955, ram_s_2_3, n2954, ram_s_2_2, 
        n2953, ram_s_2_1, n2952, n2951, ram_s_1_7, n2950, ram_s_1_6, 
        n2949, ram_s_1_5, n2948, n2947, ram_s_1_3, n2946, ram_s_1_2, 
        n2945, ram_s_1_1, n2944, n2943, ram_s_0_7, n2942, ram_s_0_6, 
        n2941, ram_s_0_5, n2940, n2939, ram_s_0_3, n2938, ram_s_0_2, 
        n2937, ram_s_0_1, n2936, n11471, n11474, n11435, n11438, 
        n8826, n8827, n11345, n8809, n8808, n11348, n9657, n9658, 
        n11339, n9280, n9279, n11342, n11264, n8806, n11315, n8800, 
        n11303, n11306, n11273, n11276, n11073, n11074, n11261, 
        n11065, n11064, n34, n6, n26, n27, n32, n7, n24, n25, 
        n30, n22, n23, n8821, n8822, n11552, n14786, n13748, 
        n11654, n12200, n14378, n12374, n12206, n12548, n28, n20, 
        n21, n29, n35, n33, n31, n12815, n10823, n12725, n12728, 
        n11879, n8867, n11549, n8846, n11861, n11864, n12683, 
        n11843, n11657, n11831, n11834, n10643, n10733, n11651, 
        n10466, n11825, n11645, n11648, n10400, n12545, n10355, 
        n10310, n8994, n8995, n11987, n8818, n10235, n10262, n12203, 
        n11762, n10127, n11948, n8948, n12197, n13217, n13220, 
        n13223, n10033, n10032, n10290, n10291, n12467, n12431, 
        n12152, n11759, n12434, n12389, n12149, n11945, n12371, 
        n9653, n9560, n13265, n13268, n13271, n13505, n13523, 
        n13526, n13565, n13568, n13721, n13724, n13739, n13742, 
        n13745, n9845, n13751, n13835, n13838, n14015, n14069, 
        n14072, n14135, n14375, n9464, n14441, n14579, n14582, 
        n14651, n14771, n14783, n14903, n14969, n15023, n15239;
    
    SB_LUT4 instruction_9__bdd_4_lut_10185 (.I0(\instruction[9] ), .I1(n11037), 
            .I2(n11038), .I3(\instruction[10] ), .O(n11231));
    defparam instruction_9__bdd_4_lut_10185.LUT_INIT = 16'he4aa;
    SB_LUT4 n11231_bdd_4_lut (.I0(n11231), .I1(n11026), .I2(n11025), .I3(\instruction[10] ), 
            .O(n11234));
    defparam n11231_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11119 (.I0(\instruction[8] ), .I1(ram_s_26_6), 
            .I2(ram_s_27_6), .I3(\instruction[9] ), .O(n12365));
    defparam instruction_8__bdd_4_lut_11119.LUT_INIT = 16'he4aa;
    SB_LUT4 instruction_8__bdd_4_lut_10501 (.I0(\instruction[8] ), .I1(ram_s_2_4), 
            .I2(ram_s_3_4), .I3(\instruction[9] ), .O(n11519));
    defparam instruction_8__bdd_4_lut_10501.LUT_INIT = 16'he4aa;
    SB_LUT4 n12365_bdd_4_lut (.I0(n12365), .I1(ram_s_25_6), .I2(ram_s_24_6), 
            .I3(\instruction[9] ), .O(n12368));
    defparam n12365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11519_bdd_4_lut (.I0(n11519), .I1(ram_s_1_4), .I2(ram_s_0_4), 
            .I3(\instruction[9] ), .O(n11522));
    defparam n11519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11808 (.I0(\instruction[8] ), .I1(ram_s_10_2), 
            .I2(ram_s_11_2), .I3(\instruction[9] ), .O(n13037));
    defparam instruction_8__bdd_4_lut_11808.LUT_INIT = 16'he4aa;
    SB_LUT4 instruction_8__bdd_4_lut_10920 (.I0(\instruction[8] ), .I1(ram_s_30_3), 
            .I2(ram_s_31_3), .I3(\instruction[9] ), .O(n12131));
    defparam instruction_8__bdd_4_lut_10920.LUT_INIT = 16'he4aa;
    SB_LUT4 n13037_bdd_4_lut (.I0(n13037), .I1(ram_s_9_2), .I2(ram_s_8_2), 
            .I3(\instruction[9] ), .O(n13040));
    defparam n13037_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12131_bdd_4_lut (.I0(n12131), .I1(ram_s_29_3), .I2(ram_s_28_3), 
            .I3(\instruction[9] ), .O(n12134));
    defparam n12131_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10750 (.I0(\instruction[8] ), .I1(ram_s_30_0), 
            .I2(ram_s_31_0), .I3(\instruction[9] ), .O(n11927));
    defparam instruction_8__bdd_4_lut_10750.LUT_INIT = 16'he4aa;
    SB_LUT4 n11927_bdd_4_lut (.I0(n11927), .I1(ram_s_29_0), .I2(ram_s_28_0), 
            .I3(\instruction[9] ), .O(n11012));
    defparam n11927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i779_780 (.Q(ram_s_31_7), .C(CLK_3P3_MHZ_c), .D(n3192));   // src/ram.vhd(56[12:17])
    SB_DFF i776_777 (.Q(ram_s_31_6), .C(CLK_3P3_MHZ_c), .D(n3191));   // src/ram.vhd(56[12:17])
    SB_LUT4 instruction_8__bdd_4_lut_10596 (.I0(\instruction[8] ), .I1(ram_s_18_0), 
            .I2(ram_s_19_0), .I3(\instruction[9] ), .O(n11741));
    defparam instruction_8__bdd_4_lut_10596.LUT_INIT = 16'he4aa;
    SB_LUT4 n11741_bdd_4_lut (.I0(n11741), .I1(ram_s_17_0), .I2(ram_s_16_0), 
            .I3(\instruction[9] ), .O(n11744));
    defparam n11741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i773_774 (.Q(ram_s_31_5), .C(CLK_3P3_MHZ_c), .D(n3190));   // src/ram.vhd(56[12:17])
    SB_DFF i770_771 (.Q(ram_s_31_4), .C(CLK_3P3_MHZ_c), .D(n3189));   // src/ram.vhd(56[12:17])
    SB_DFF i767_768 (.Q(ram_s_31_3), .C(CLK_3P3_MHZ_c), .D(n3188));   // src/ram.vhd(56[12:17])
    SB_DFF i764_765 (.Q(ram_s_31_2), .C(CLK_3P3_MHZ_c), .D(n3187));   // src/ram.vhd(56[12:17])
    SB_DFF i761_762 (.Q(ram_s_31_1), .C(CLK_3P3_MHZ_c), .D(n3186));   // src/ram.vhd(56[12:17])
    SB_DFF i758_759 (.Q(ram_s_31_0), .C(CLK_3P3_MHZ_c), .D(n3185));   // src/ram.vhd(56[12:17])
    SB_LUT4 instruction_10__bdd_4_lut_10960 (.I0(\instruction[10] ), .I1(n11846), 
            .I2(n11828), .I3(\instruction[11] ), .O(n11915));
    defparam instruction_10__bdd_4_lut_10960.LUT_INIT = 16'he4aa;
    SB_LUT4 n11915_bdd_4_lut (.I0(n11915), .I1(n11882), .I2(n11900), .I3(\instruction[11] ), 
            .O(n11918));
    defparam n11915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10905 (.I0(\instruction[8] ), .I1(ram_s_26_2), 
            .I2(ram_s_27_2), .I3(\instruction[9] ), .O(n12101));
    defparam instruction_8__bdd_4_lut_10905.LUT_INIT = 16'he4aa;
    SB_LUT4 instruction_8__bdd_4_lut_11658 (.I0(\instruction[8] ), .I1(ram_s_30_7), 
            .I2(ram_s_31_7), .I3(\instruction[9] ), .O(n12995));
    defparam instruction_8__bdd_4_lut_11658.LUT_INIT = 16'he4aa;
    SB_DFF i755_756 (.Q(ram_s_30_7), .C(CLK_3P3_MHZ_c), .D(n3184));   // src/ram.vhd(56[12:17])
    SB_DFF i752_753 (.Q(ram_s_30_6), .C(CLK_3P3_MHZ_c), .D(n3183));   // src/ram.vhd(56[12:17])
    SB_DFF i749_750 (.Q(ram_s_30_5), .C(CLK_3P3_MHZ_c), .D(n3182));   // src/ram.vhd(56[12:17])
    SB_DFF i746_747 (.Q(ram_s_30_4), .C(CLK_3P3_MHZ_c), .D(n3181));   // src/ram.vhd(56[12:17])
    SB_LUT4 n12995_bdd_4_lut (.I0(n12995), .I1(ram_s_29_7), .I2(ram_s_28_7), 
            .I3(\instruction[9] ), .O(n10421));
    defparam n12995_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12101_bdd_4_lut (.I0(n12101), .I1(ram_s_25_2), .I2(ram_s_24_2), 
            .I3(\instruction[9] ), .O(n8858));
    defparam n12101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i743_744 (.Q(ram_s_30_3), .C(CLK_3P3_MHZ_c), .D(n3180));   // src/ram.vhd(56[12:17])
    SB_LUT4 instruction_8__bdd_4_lut_11623 (.I0(\instruction[8] ), .I1(ram_s_14_2), 
            .I2(ram_s_15_2), .I3(\instruction[9] ), .O(n12977));
    defparam instruction_8__bdd_4_lut_11623.LUT_INIT = 16'he4aa;
    SB_LUT4 n12977_bdd_4_lut (.I0(n12977), .I1(ram_s_13_2), .I2(ram_s_12_2), 
            .I3(\instruction[9] ), .O(n12980));
    defparam n12977_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i740_741 (.Q(ram_s_30_2), .C(CLK_3P3_MHZ_c), .D(n3179));   // src/ram.vhd(56[12:17])
    SB_DFF i737_738 (.Q(ram_s_30_1), .C(CLK_3P3_MHZ_c), .D(n3178));   // src/ram.vhd(56[12:17])
    SB_DFF i734_735 (.Q(ram_s_30_0), .C(CLK_3P3_MHZ_c), .D(n3177));   // src/ram.vhd(56[12:17])
    SB_DFF i731_732 (.Q(ram_s_29_7), .C(CLK_3P3_MHZ_c), .D(n3176));   // src/ram.vhd(56[12:17])
    SB_DFF i728_729 (.Q(ram_s_29_6), .C(CLK_3P3_MHZ_c), .D(n3174));   // src/ram.vhd(56[12:17])
    SB_DFF i725_726 (.Q(ram_s_29_5), .C(CLK_3P3_MHZ_c), .D(n3173));   // src/ram.vhd(56[12:17])
    SB_DFF i722_723 (.Q(ram_s_29_4), .C(CLK_3P3_MHZ_c), .D(n3172));   // src/ram.vhd(56[12:17])
    SB_DFF i719_720 (.Q(ram_s_29_3), .C(CLK_3P3_MHZ_c), .D(n3171));   // src/ram.vhd(56[12:17])
    SB_DFF i716_717 (.Q(ram_s_29_2), .C(CLK_3P3_MHZ_c), .D(n3170));   // src/ram.vhd(56[12:17])
    SB_DFF i713_714 (.Q(ram_s_29_1), .C(CLK_3P3_MHZ_c), .D(n3169));   // src/ram.vhd(56[12:17])
    SB_DFF i710_711 (.Q(ram_s_29_0), .C(CLK_3P3_MHZ_c), .D(n3168));   // src/ram.vhd(56[12:17])
    SB_LUT4 instruction_10__bdd_4_lut_10725 (.I0(\instruction[10] ), .I1(n11492), 
            .I2(n11012), .I3(\instruction[11] ), .O(n11903));
    defparam instruction_10__bdd_4_lut_10725.LUT_INIT = 16'he4aa;
    SB_DFF i707_708 (.Q(ram_s_28_7), .C(CLK_3P3_MHZ_c), .D(n3167));   // src/ram.vhd(56[12:17])
    SB_LUT4 n11903_bdd_4_lut (.I0(n11903), .I1(n11498), .I2(n11744), .I3(\instruction[11] ), 
            .O(n11906));
    defparam n11903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i704_705 (.Q(ram_s_28_6), .C(CLK_3P3_MHZ_c), .D(n3166));   // src/ram.vhd(56[12:17])
    SB_DFF i701_702 (.Q(ram_s_28_5), .C(CLK_3P3_MHZ_c), .D(n3165));   // src/ram.vhd(56[12:17])
    SB_DFF i698_699 (.Q(ram_s_28_4), .C(CLK_3P3_MHZ_c), .D(n3164));   // src/ram.vhd(56[12:17])
    SB_DFF i695_696 (.Q(ram_s_28_3), .C(CLK_3P3_MHZ_c), .D(n3163));   // src/ram.vhd(56[12:17])
    SB_DFF i692_693 (.Q(ram_s_28_2), .C(CLK_3P3_MHZ_c), .D(n3162));   // src/ram.vhd(56[12:17])
    SB_DFF i689_690 (.Q(ram_s_28_1), .C(CLK_3P3_MHZ_c), .D(n3161));   // src/ram.vhd(56[12:17])
    SB_DFF i686_687 (.Q(ram_s_28_0), .C(CLK_3P3_MHZ_c), .D(n3160));   // src/ram.vhd(56[12:17])
    SB_DFF i683_684 (.Q(ram_s_27_7), .C(CLK_3P3_MHZ_c), .D(n3159));   // src/ram.vhd(56[12:17])
    SB_DFF i680_681 (.Q(ram_s_27_6), .C(CLK_3P3_MHZ_c), .D(n3158));   // src/ram.vhd(56[12:17])
    SB_DFF i677_678 (.Q(ram_s_27_5), .C(CLK_3P3_MHZ_c), .D(n3157));   // src/ram.vhd(56[12:17])
    SB_DFF i674_675 (.Q(ram_s_27_4), .C(CLK_3P3_MHZ_c), .D(n3156));   // src/ram.vhd(56[12:17])
    SB_DFF i671_672 (.Q(ram_s_27_3), .C(CLK_3P3_MHZ_c), .D(n3155));   // src/ram.vhd(56[12:17])
    SB_DFF i668_669 (.Q(ram_s_27_2), .C(CLK_3P3_MHZ_c), .D(n3154));   // src/ram.vhd(56[12:17])
    SB_DFF i665_666 (.Q(ram_s_27_1), .C(CLK_3P3_MHZ_c), .D(n3153));   // src/ram.vhd(56[12:17])
    SB_DFF i662_663 (.Q(ram_s_27_0), .C(CLK_3P3_MHZ_c), .D(n3152));   // src/ram.vhd(56[12:17])
    SB_DFF i659_660 (.Q(ram_s_26_7), .C(CLK_3P3_MHZ_c), .D(n3151));   // src/ram.vhd(56[12:17])
    SB_DFF i656_657 (.Q(ram_s_26_6), .C(CLK_3P3_MHZ_c), .D(n3150));   // src/ram.vhd(56[12:17])
    SB_DFF i653_654 (.Q(ram_s_26_5), .C(CLK_3P3_MHZ_c), .D(n3149));   // src/ram.vhd(56[12:17])
    SB_DFF i650_651 (.Q(ram_s_26_4), .C(CLK_3P3_MHZ_c), .D(n3148));   // src/ram.vhd(56[12:17])
    SB_DFF i647_648 (.Q(ram_s_26_3), .C(CLK_3P3_MHZ_c), .D(n3147));   // src/ram.vhd(56[12:17])
    SB_DFF i644_645 (.Q(ram_s_26_2), .C(CLK_3P3_MHZ_c), .D(n3146));   // src/ram.vhd(56[12:17])
    SB_DFF i641_642 (.Q(ram_s_26_1), .C(CLK_3P3_MHZ_c), .D(n3145));   // src/ram.vhd(56[12:17])
    SB_DFF i638_639 (.Q(ram_s_26_0), .C(CLK_3P3_MHZ_c), .D(n3144));   // src/ram.vhd(56[12:17])
    SB_DFF i635_636 (.Q(ram_s_25_7), .C(CLK_3P3_MHZ_c), .D(n3143));   // src/ram.vhd(56[12:17])
    SB_DFF i632_633 (.Q(ram_s_25_6), .C(CLK_3P3_MHZ_c), .D(n3142));   // src/ram.vhd(56[12:17])
    SB_DFF i629_630 (.Q(ram_s_25_5), .C(CLK_3P3_MHZ_c), .D(n3141));   // src/ram.vhd(56[12:17])
    SB_DFF i626_627 (.Q(ram_s_25_4), .C(CLK_3P3_MHZ_c), .D(n3140));   // src/ram.vhd(56[12:17])
    SB_DFF i623_624 (.Q(ram_s_25_3), .C(CLK_3P3_MHZ_c), .D(n3139));   // src/ram.vhd(56[12:17])
    SB_DFF i620_621 (.Q(ram_s_25_2), .C(CLK_3P3_MHZ_c), .D(n3138));   // src/ram.vhd(56[12:17])
    SB_DFF i617_618 (.Q(ram_s_25_1), .C(CLK_3P3_MHZ_c), .D(n3137));   // src/ram.vhd(56[12:17])
    SB_DFF i614_615 (.Q(ram_s_25_0), .C(CLK_3P3_MHZ_c), .D(n3136));   // src/ram.vhd(56[12:17])
    SB_DFF i611_612 (.Q(ram_s_24_7), .C(CLK_3P3_MHZ_c), .D(n3135));   // src/ram.vhd(56[12:17])
    SB_DFF i608_609 (.Q(ram_s_24_6), .C(CLK_3P3_MHZ_c), .D(n3134));   // src/ram.vhd(56[12:17])
    SB_DFF i605_606 (.Q(ram_s_24_5), .C(CLK_3P3_MHZ_c), .D(n3133));   // src/ram.vhd(56[12:17])
    SB_DFF i602_603 (.Q(ram_s_24_4), .C(CLK_3P3_MHZ_c), .D(n3132));   // src/ram.vhd(56[12:17])
    SB_DFF i599_600 (.Q(ram_s_24_3), .C(CLK_3P3_MHZ_c), .D(n3131));   // src/ram.vhd(56[12:17])
    SB_DFF i596_597 (.Q(ram_s_24_2), .C(CLK_3P3_MHZ_c), .D(n3130));   // src/ram.vhd(56[12:17])
    SB_DFF i593_594 (.Q(ram_s_24_1), .C(CLK_3P3_MHZ_c), .D(n3129));   // src/ram.vhd(56[12:17])
    SB_DFF i590_591 (.Q(ram_s_24_0), .C(CLK_3P3_MHZ_c), .D(n3128));   // src/ram.vhd(56[12:17])
    SB_DFF i587_588 (.Q(ram_s_23_7), .C(CLK_3P3_MHZ_c), .D(n3127));   // src/ram.vhd(56[12:17])
    SB_DFF i584_585 (.Q(ram_s_23_6), .C(CLK_3P3_MHZ_c), .D(n3126));   // src/ram.vhd(56[12:17])
    SB_DFF i581_582 (.Q(ram_s_23_5), .C(CLK_3P3_MHZ_c), .D(n3125));   // src/ram.vhd(56[12:17])
    SB_LUT4 instruction_8__bdd_4_lut_10397 (.I0(\instruction[8] ), .I1(ram_s_22_0), 
            .I2(ram_s_23_0), .I3(\instruction[9] ), .O(n11495));
    defparam instruction_8__bdd_4_lut_10397.LUT_INIT = 16'he4aa;
    SB_LUT4 instruction_8__bdd_4_lut_10735 (.I0(\instruction[8] ), .I1(ram_s_2_0), 
            .I2(ram_s_3_0), .I3(\instruction[9] ), .O(n11897));
    defparam instruction_8__bdd_4_lut_10735.LUT_INIT = 16'he4aa;
    SB_LUT4 n11495_bdd_4_lut (.I0(n11495), .I1(ram_s_21_0), .I2(ram_s_20_0), 
            .I3(\instruction[9] ), .O(n11498));
    defparam n11495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i578_579 (.Q(ram_s_23_4), .C(CLK_3P3_MHZ_c), .D(n3124));   // src/ram.vhd(56[12:17])
    SB_DFF i575_576 (.Q(ram_s_23_3), .C(CLK_3P3_MHZ_c), .D(n3123));   // src/ram.vhd(56[12:17])
    SB_DFF i572_573 (.Q(ram_s_23_2), .C(CLK_3P3_MHZ_c), .D(n3122));   // src/ram.vhd(56[12:17])
    SB_DFF i569_570 (.Q(ram_s_23_1), .C(CLK_3P3_MHZ_c), .D(n3121));   // src/ram.vhd(56[12:17])
    SB_DFF i566_567 (.Q(ram_s_23_0), .C(CLK_3P3_MHZ_c), .D(n3120));   // src/ram.vhd(56[12:17])
    SB_DFF i563_564 (.Q(ram_s_22_7), .C(CLK_3P3_MHZ_c), .D(n3119));   // src/ram.vhd(56[12:17])
    SB_DFF i560_561 (.Q(ram_s_22_6), .C(CLK_3P3_MHZ_c), .D(n3118));   // src/ram.vhd(56[12:17])
    SB_DFF i557_558 (.Q(ram_s_22_5), .C(CLK_3P3_MHZ_c), .D(n3117));   // src/ram.vhd(56[12:17])
    SB_DFF i554_555 (.Q(ram_s_22_4), .C(CLK_3P3_MHZ_c), .D(n3116));   // src/ram.vhd(56[12:17])
    SB_LUT4 n11897_bdd_4_lut (.I0(n11897), .I1(ram_s_1_0), .I2(ram_s_0_0), 
            .I3(\instruction[9] ), .O(n11900));
    defparam n11897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10377 (.I0(\instruction[8] ), .I1(ram_s_26_0), 
            .I2(ram_s_27_0), .I3(\instruction[9] ), .O(n11489));
    defparam instruction_8__bdd_4_lut_10377.LUT_INIT = 16'he4aa;
    SB_DFF i551_552 (.Q(ram_s_22_3), .C(CLK_3P3_MHZ_c), .D(n3115));   // src/ram.vhd(56[12:17])
    SB_DFF i548_549 (.Q(ram_s_22_2), .C(CLK_3P3_MHZ_c), .D(n3114));   // src/ram.vhd(56[12:17])
    SB_DFF i545_546 (.Q(ram_s_22_1), .C(CLK_3P3_MHZ_c), .D(n3113));   // src/ram.vhd(56[12:17])
    SB_DFF i542_543 (.Q(ram_s_22_0), .C(CLK_3P3_MHZ_c), .D(n3112));   // src/ram.vhd(56[12:17])
    SB_DFF i539_540 (.Q(ram_s_21_7), .C(CLK_3P3_MHZ_c), .D(n3111));   // src/ram.vhd(56[12:17])
    SB_DFF i536_537 (.Q(ram_s_21_6), .C(CLK_3P3_MHZ_c), .D(n3110));   // src/ram.vhd(56[12:17])
    SB_DFF i533_534 (.Q(ram_s_21_5), .C(CLK_3P3_MHZ_c), .D(n3109));   // src/ram.vhd(56[12:17])
    SB_DFF i530_531 (.Q(ram_s_21_4), .C(CLK_3P3_MHZ_c), .D(n3108));   // src/ram.vhd(56[12:17])
    SB_LUT4 instruction_8__bdd_4_lut_11608 (.I0(\instruction[8] ), .I1(ram_s_18_2), 
            .I2(ram_s_19_2), .I3(\instruction[9] ), .O(n12923));
    defparam instruction_8__bdd_4_lut_11608.LUT_INIT = 16'he4aa;
    SB_DFF i527_528 (.Q(ram_s_21_3), .C(CLK_3P3_MHZ_c), .D(n3107));   // src/ram.vhd(56[12:17])
    SB_DFF i524_525 (.Q(ram_s_21_2), .C(CLK_3P3_MHZ_c), .D(n3106));   // src/ram.vhd(56[12:17])
    SB_DFF i521_522 (.Q(ram_s_21_1), .C(CLK_3P3_MHZ_c), .D(n3105));   // src/ram.vhd(56[12:17])
    SB_DFF i518_519 (.Q(ram_s_21_0), .C(CLK_3P3_MHZ_c), .D(n3104));   // src/ram.vhd(56[12:17])
    SB_DFF i515_516 (.Q(ram_s_20_7), .C(CLK_3P3_MHZ_c), .D(n3103));   // src/ram.vhd(56[12:17])
    SB_DFF i512_513 (.Q(ram_s_20_6), .C(CLK_3P3_MHZ_c), .D(n3102));   // src/ram.vhd(56[12:17])
    SB_DFF i509_510 (.Q(ram_s_20_5), .C(CLK_3P3_MHZ_c), .D(n3101));   // src/ram.vhd(56[12:17])
    SB_DFF i506_507 (.Q(ram_s_20_4), .C(CLK_3P3_MHZ_c), .D(n3100));   // src/ram.vhd(56[12:17])
    SB_DFF i503_504 (.Q(ram_s_20_3), .C(CLK_3P3_MHZ_c), .D(n3099));   // src/ram.vhd(56[12:17])
    SB_DFF i500_501 (.Q(ram_s_20_2), .C(CLK_3P3_MHZ_c), .D(n3098));   // src/ram.vhd(56[12:17])
    SB_DFF i497_498 (.Q(ram_s_20_1), .C(CLK_3P3_MHZ_c), .D(n3097));   // src/ram.vhd(56[12:17])
    SB_DFF i494_495 (.Q(ram_s_20_0), .C(CLK_3P3_MHZ_c), .D(n3096));   // src/ram.vhd(56[12:17])
    SB_DFF i491_492 (.Q(ram_s_19_7), .C(CLK_3P3_MHZ_c), .D(n3095));   // src/ram.vhd(56[12:17])
    SB_DFF i488_489 (.Q(ram_s_19_6), .C(CLK_3P3_MHZ_c), .D(n3094));   // src/ram.vhd(56[12:17])
    SB_DFF i485_486 (.Q(ram_s_19_5), .C(CLK_3P3_MHZ_c), .D(n3093));   // src/ram.vhd(56[12:17])
    SB_DFF i482_483 (.Q(ram_s_19_4), .C(CLK_3P3_MHZ_c), .D(n3092));   // src/ram.vhd(56[12:17])
    SB_DFF i479_480 (.Q(ram_s_19_3), .C(CLK_3P3_MHZ_c), .D(n3091));   // src/ram.vhd(56[12:17])
    SB_DFF i476_477 (.Q(ram_s_19_2), .C(CLK_3P3_MHZ_c), .D(n3090));   // src/ram.vhd(56[12:17])
    SB_DFF i473_474 (.Q(ram_s_19_1), .C(CLK_3P3_MHZ_c), .D(n3089));   // src/ram.vhd(56[12:17])
    SB_DFF i470_471 (.Q(ram_s_19_0), .C(CLK_3P3_MHZ_c), .D(n3088));   // src/ram.vhd(56[12:17])
    SB_DFF i467_468 (.Q(ram_s_18_7), .C(CLK_3P3_MHZ_c), .D(n3087));   // src/ram.vhd(56[12:17])
    SB_DFF i464_465 (.Q(ram_s_18_6), .C(CLK_3P3_MHZ_c), .D(n3086));   // src/ram.vhd(56[12:17])
    SB_DFF i461_462 (.Q(ram_s_18_5), .C(CLK_3P3_MHZ_c), .D(n3085));   // src/ram.vhd(56[12:17])
    SB_LUT4 n12923_bdd_4_lut (.I0(n12923), .I1(ram_s_17_2), .I2(ram_s_16_2), 
            .I3(\instruction[9] ), .O(n8840));
    defparam n12923_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i458_459 (.Q(ram_s_18_4), .C(CLK_3P3_MHZ_c), .D(n3084));   // src/ram.vhd(56[12:17])
    SB_DFF i455_456 (.Q(ram_s_18_3), .C(CLK_3P3_MHZ_c), .D(n3083));   // src/ram.vhd(56[12:17])
    SB_DFF i452_453 (.Q(ram_s_18_2), .C(CLK_3P3_MHZ_c), .D(n3082));   // src/ram.vhd(56[12:17])
    SB_DFF i449_450 (.Q(ram_s_18_1), .C(CLK_3P3_MHZ_c), .D(n3081));   // src/ram.vhd(56[12:17])
    SB_DFF i446_447 (.Q(ram_s_18_0), .C(CLK_3P3_MHZ_c), .D(n3080));   // src/ram.vhd(56[12:17])
    SB_DFF i443_444 (.Q(ram_s_17_7), .C(CLK_3P3_MHZ_c), .D(n3079));   // src/ram.vhd(56[12:17])
    SB_DFF i440_441 (.Q(ram_s_17_6), .C(CLK_3P3_MHZ_c), .D(n3078));   // src/ram.vhd(56[12:17])
    SB_DFF i437_438 (.Q(ram_s_17_5), .C(CLK_3P3_MHZ_c), .D(n3077));   // src/ram.vhd(56[12:17])
    SB_DFF i434_435 (.Q(ram_s_17_4), .C(CLK_3P3_MHZ_c), .D(n3076));   // src/ram.vhd(56[12:17])
    SB_DFF i431_432 (.Q(ram_s_17_3), .C(CLK_3P3_MHZ_c), .D(n3075));   // src/ram.vhd(56[12:17])
    SB_DFF i428_429 (.Q(ram_s_17_2), .C(CLK_3P3_MHZ_c), .D(n3074));   // src/ram.vhd(56[12:17])
    SB_DFF i425_426 (.Q(ram_s_17_1), .C(CLK_3P3_MHZ_c), .D(n3073));   // src/ram.vhd(56[12:17])
    SB_LUT4 n11489_bdd_4_lut (.I0(n11489), .I1(ram_s_25_0), .I2(ram_s_24_0), 
            .I3(\instruction[9] ), .O(n11492));
    defparam n11489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i422_423 (.Q(ram_s_17_0), .C(CLK_3P3_MHZ_c), .D(n3072));   // src/ram.vhd(56[12:17])
    SB_DFF i419_420 (.Q(ram_s_16_7), .C(CLK_3P3_MHZ_c), .D(n3071));   // src/ram.vhd(56[12:17])
    SB_DFF i416_417 (.Q(ram_s_16_6), .C(CLK_3P3_MHZ_c), .D(n3070));   // src/ram.vhd(56[12:17])
    SB_DFF i413_414 (.Q(ram_s_16_5), .C(CLK_3P3_MHZ_c), .D(n3069));   // src/ram.vhd(56[12:17])
    SB_DFF i410_411 (.Q(ram_s_16_4), .C(CLK_3P3_MHZ_c), .D(n3068));   // src/ram.vhd(56[12:17])
    SB_DFF i407_408 (.Q(ram_s_16_3), .C(CLK_3P3_MHZ_c), .D(n3067));   // src/ram.vhd(56[12:17])
    SB_DFF i404_405 (.Q(ram_s_16_2), .C(CLK_3P3_MHZ_c), .D(n3066));   // src/ram.vhd(56[12:17])
    SB_DFF i401_402 (.Q(ram_s_16_1), .C(CLK_3P3_MHZ_c), .D(n3065));   // src/ram.vhd(56[12:17])
    SB_DFF i398_399 (.Q(ram_s_16_0), .C(CLK_3P3_MHZ_c), .D(n3064));   // src/ram.vhd(56[12:17])
    SB_DFF i395_396 (.Q(ram_s_15_7), .C(CLK_3P3_MHZ_c), .D(n3063));   // src/ram.vhd(56[12:17])
    SB_DFF i392_393 (.Q(ram_s_15_6), .C(CLK_3P3_MHZ_c), .D(n3062));   // src/ram.vhd(56[12:17])
    SB_DFF i389_390 (.Q(ram_s_15_5), .C(CLK_3P3_MHZ_c), .D(n3061));   // src/ram.vhd(56[12:17])
    SB_DFF i386_387 (.Q(ram_s_15_4), .C(CLK_3P3_MHZ_c), .D(n3060));   // src/ram.vhd(56[12:17])
    SB_DFF i383_384 (.Q(ram_s_15_3), .C(CLK_3P3_MHZ_c), .D(n3059));   // src/ram.vhd(56[12:17])
    SB_DFF i380_381 (.Q(ram_s_15_2), .C(CLK_3P3_MHZ_c), .D(n3058));   // src/ram.vhd(56[12:17])
    SB_DFF i377_378 (.Q(ram_s_15_1), .C(CLK_3P3_MHZ_c), .D(n3057));   // src/ram.vhd(56[12:17])
    SB_DFF i374_375 (.Q(ram_s_15_0), .C(CLK_3P3_MHZ_c), .D(n3056));   // src/ram.vhd(56[12:17])
    SB_DFF i371_372 (.Q(ram_s_14_7), .C(CLK_3P3_MHZ_c), .D(n3055));   // src/ram.vhd(56[12:17])
    SB_DFF i368_369 (.Q(ram_s_14_6), .C(CLK_3P3_MHZ_c), .D(n3054));   // src/ram.vhd(56[12:17])
    SB_DFF i365_366 (.Q(ram_s_14_5), .C(CLK_3P3_MHZ_c), .D(n3053));   // src/ram.vhd(56[12:17])
    SB_DFF i362_363 (.Q(ram_s_14_4), .C(CLK_3P3_MHZ_c), .D(n3052));   // src/ram.vhd(56[12:17])
    SB_DFF i359_360 (.Q(ram_s_14_3), .C(CLK_3P3_MHZ_c), .D(n3051));   // src/ram.vhd(56[12:17])
    SB_DFF i356_357 (.Q(ram_s_14_2), .C(CLK_3P3_MHZ_c), .D(n3050));   // src/ram.vhd(56[12:17])
    SB_DFF i353_354 (.Q(ram_s_14_1), .C(CLK_3P3_MHZ_c), .D(n3049));   // src/ram.vhd(56[12:17])
    SB_DFF i350_351 (.Q(ram_s_14_0), .C(CLK_3P3_MHZ_c), .D(n3048));   // src/ram.vhd(56[12:17])
    SB_DFF i347_348 (.Q(ram_s_13_7), .C(CLK_3P3_MHZ_c), .D(n3047));   // src/ram.vhd(56[12:17])
    SB_DFF i344_345 (.Q(ram_s_13_6), .C(CLK_3P3_MHZ_c), .D(n3046));   // src/ram.vhd(56[12:17])
    SB_DFF i341_342 (.Q(ram_s_13_5), .C(CLK_3P3_MHZ_c), .D(n3045));   // src/ram.vhd(56[12:17])
    SB_DFF i338_339 (.Q(ram_s_13_4), .C(CLK_3P3_MHZ_c), .D(n3044));   // src/ram.vhd(56[12:17])
    SB_DFF i335_336 (.Q(ram_s_13_3), .C(CLK_3P3_MHZ_c), .D(n3043));   // src/ram.vhd(56[12:17])
    SB_DFF i332_333 (.Q(ram_s_13_2), .C(CLK_3P3_MHZ_c), .D(n3042));   // src/ram.vhd(56[12:17])
    SB_DFF i329_330 (.Q(ram_s_13_1), .C(CLK_3P3_MHZ_c), .D(n3041));   // src/ram.vhd(56[12:17])
    SB_DFF i326_327 (.Q(ram_s_13_0), .C(CLK_3P3_MHZ_c), .D(n3040));   // src/ram.vhd(56[12:17])
    SB_DFF i323_324 (.Q(ram_s_12_7), .C(CLK_3P3_MHZ_c), .D(n3039));   // src/ram.vhd(56[12:17])
    SB_DFF i320_321 (.Q(ram_s_12_6), .C(CLK_3P3_MHZ_c), .D(n3038));   // src/ram.vhd(56[12:17])
    SB_DFF i317_318 (.Q(ram_s_12_5), .C(CLK_3P3_MHZ_c), .D(n3037));   // src/ram.vhd(56[12:17])
    SB_DFF i314_315 (.Q(ram_s_12_4), .C(CLK_3P3_MHZ_c), .D(n3036));   // src/ram.vhd(56[12:17])
    SB_DFF i311_312 (.Q(ram_s_12_3), .C(CLK_3P3_MHZ_c), .D(n3035));   // src/ram.vhd(56[12:17])
    SB_DFF i308_309 (.Q(ram_s_12_2), .C(CLK_3P3_MHZ_c), .D(n3034));   // src/ram.vhd(56[12:17])
    SB_DFF i305_306 (.Q(ram_s_12_1), .C(CLK_3P3_MHZ_c), .D(n3033));   // src/ram.vhd(56[12:17])
    SB_DFF i302_303 (.Q(ram_s_12_0), .C(CLK_3P3_MHZ_c), .D(n3032));   // src/ram.vhd(56[12:17])
    SB_DFF i299_300 (.Q(ram_s_11_7), .C(CLK_3P3_MHZ_c), .D(n3031));   // src/ram.vhd(56[12:17])
    SB_DFF i296_297 (.Q(ram_s_11_6), .C(CLK_3P3_MHZ_c), .D(n3030));   // src/ram.vhd(56[12:17])
    SB_DFF i293_294 (.Q(ram_s_11_5), .C(CLK_3P3_MHZ_c), .D(n3029));   // src/ram.vhd(56[12:17])
    SB_DFF i290_291 (.Q(ram_s_11_4), .C(CLK_3P3_MHZ_c), .D(n3028));   // src/ram.vhd(56[12:17])
    SB_DFF i287_288 (.Q(ram_s_11_3), .C(CLK_3P3_MHZ_c), .D(n3027));   // src/ram.vhd(56[12:17])
    SB_DFF i284_285 (.Q(ram_s_11_2), .C(CLK_3P3_MHZ_c), .D(n3026));   // src/ram.vhd(56[12:17])
    SB_DFF i281_282 (.Q(ram_s_11_1), .C(CLK_3P3_MHZ_c), .D(n3025));   // src/ram.vhd(56[12:17])
    SB_DFF i278_279 (.Q(ram_s_11_0), .C(CLK_3P3_MHZ_c), .D(n3024));   // src/ram.vhd(56[12:17])
    SB_DFF i275_276 (.Q(ram_s_10_7), .C(CLK_3P3_MHZ_c), .D(n3023));   // src/ram.vhd(56[12:17])
    SB_DFF i272_273 (.Q(ram_s_10_6), .C(CLK_3P3_MHZ_c), .D(n3022));   // src/ram.vhd(56[12:17])
    SB_DFF i269_270 (.Q(ram_s_10_5), .C(CLK_3P3_MHZ_c), .D(n3021));   // src/ram.vhd(56[12:17])
    SB_DFF i266_267 (.Q(ram_s_10_4), .C(CLK_3P3_MHZ_c), .D(n3020));   // src/ram.vhd(56[12:17])
    SB_DFF i263_264 (.Q(ram_s_10_3), .C(CLK_3P3_MHZ_c), .D(n3019));   // src/ram.vhd(56[12:17])
    SB_DFF i260_261 (.Q(ram_s_10_2), .C(CLK_3P3_MHZ_c), .D(n3018));   // src/ram.vhd(56[12:17])
    SB_DFF i257_258 (.Q(ram_s_10_1), .C(CLK_3P3_MHZ_c), .D(n3017));   // src/ram.vhd(56[12:17])
    SB_DFF i254_255 (.Q(ram_s_10_0), .C(CLK_3P3_MHZ_c), .D(n3016));   // src/ram.vhd(56[12:17])
    SB_DFF i251_252 (.Q(ram_s_9_7), .C(CLK_3P3_MHZ_c), .D(n3015));   // src/ram.vhd(56[12:17])
    SB_DFF i248_249 (.Q(ram_s_9_6), .C(CLK_3P3_MHZ_c), .D(n3014));   // src/ram.vhd(56[12:17])
    SB_DFF i245_246 (.Q(ram_s_9_5), .C(CLK_3P3_MHZ_c), .D(n3013));   // src/ram.vhd(56[12:17])
    SB_DFF i242_243 (.Q(ram_s_9_4), .C(CLK_3P3_MHZ_c), .D(n3012));   // src/ram.vhd(56[12:17])
    SB_DFF i239_240 (.Q(ram_s_9_3), .C(CLK_3P3_MHZ_c), .D(n3011));   // src/ram.vhd(56[12:17])
    SB_DFF i236_237 (.Q(ram_s_9_2), .C(CLK_3P3_MHZ_c), .D(n3010));   // src/ram.vhd(56[12:17])
    SB_DFF i233_234 (.Q(ram_s_9_1), .C(CLK_3P3_MHZ_c), .D(n3009));   // src/ram.vhd(56[12:17])
    SB_DFF i230_231 (.Q(ram_s_9_0), .C(CLK_3P3_MHZ_c), .D(n3008));   // src/ram.vhd(56[12:17])
    SB_DFF i227_228 (.Q(ram_s_8_7), .C(CLK_3P3_MHZ_c), .D(n3007));   // src/ram.vhd(56[12:17])
    SB_DFF i224_225 (.Q(ram_s_8_6), .C(CLK_3P3_MHZ_c), .D(n3006));   // src/ram.vhd(56[12:17])
    SB_DFF i221_222 (.Q(ram_s_8_5), .C(CLK_3P3_MHZ_c), .D(n3005));   // src/ram.vhd(56[12:17])
    SB_DFF i218_219 (.Q(ram_s_8_4), .C(CLK_3P3_MHZ_c), .D(n3004));   // src/ram.vhd(56[12:17])
    SB_DFF i215_216 (.Q(ram_s_8_3), .C(CLK_3P3_MHZ_c), .D(n3003));   // src/ram.vhd(56[12:17])
    SB_DFF i212_213 (.Q(ram_s_8_2), .C(CLK_3P3_MHZ_c), .D(n3002));   // src/ram.vhd(56[12:17])
    SB_DFF i209_210 (.Q(ram_s_8_1), .C(CLK_3P3_MHZ_c), .D(n3001));   // src/ram.vhd(56[12:17])
    SB_DFF i206_207 (.Q(ram_s_8_0), .C(CLK_3P3_MHZ_c), .D(n3000));   // src/ram.vhd(56[12:17])
    SB_DFF i203_204 (.Q(ram_s_7_7), .C(CLK_3P3_MHZ_c), .D(n2999));   // src/ram.vhd(56[12:17])
    SB_DFF i200_201 (.Q(ram_s_7_6), .C(CLK_3P3_MHZ_c), .D(n2998));   // src/ram.vhd(56[12:17])
    SB_DFF i197_198 (.Q(ram_s_7_5), .C(CLK_3P3_MHZ_c), .D(n2997));   // src/ram.vhd(56[12:17])
    SB_DFF i194_195 (.Q(ram_s_7_4), .C(CLK_3P3_MHZ_c), .D(n2996));   // src/ram.vhd(56[12:17])
    SB_DFF i191_192 (.Q(ram_s_7_3), .C(CLK_3P3_MHZ_c), .D(n2995));   // src/ram.vhd(56[12:17])
    SB_DFF i188_189 (.Q(ram_s_7_2), .C(CLK_3P3_MHZ_c), .D(n2994));   // src/ram.vhd(56[12:17])
    SB_DFF i185_186 (.Q(ram_s_7_1), .C(CLK_3P3_MHZ_c), .D(n2993));   // src/ram.vhd(56[12:17])
    SB_DFF i182_183 (.Q(ram_s_7_0), .C(CLK_3P3_MHZ_c), .D(n2992));   // src/ram.vhd(56[12:17])
    SB_DFF i179_180 (.Q(ram_s_6_7), .C(CLK_3P3_MHZ_c), .D(n2991));   // src/ram.vhd(56[12:17])
    SB_DFF i176_177 (.Q(ram_s_6_6), .C(CLK_3P3_MHZ_c), .D(n2990));   // src/ram.vhd(56[12:17])
    SB_DFF i173_174 (.Q(ram_s_6_5), .C(CLK_3P3_MHZ_c), .D(n2989));   // src/ram.vhd(56[12:17])
    SB_DFF i170_171 (.Q(ram_s_6_4), .C(CLK_3P3_MHZ_c), .D(n2988));   // src/ram.vhd(56[12:17])
    SB_DFF i167_168 (.Q(ram_s_6_3), .C(CLK_3P3_MHZ_c), .D(n2987));   // src/ram.vhd(56[12:17])
    SB_DFF i164_165 (.Q(ram_s_6_2), .C(CLK_3P3_MHZ_c), .D(n2986));   // src/ram.vhd(56[12:17])
    SB_DFF i161_162 (.Q(ram_s_6_1), .C(CLK_3P3_MHZ_c), .D(n2985));   // src/ram.vhd(56[12:17])
    SB_DFF i158_159 (.Q(ram_s_6_0), .C(CLK_3P3_MHZ_c), .D(n2984));   // src/ram.vhd(56[12:17])
    SB_DFF i155_156 (.Q(ram_s_5_7), .C(CLK_3P3_MHZ_c), .D(n2983));   // src/ram.vhd(56[12:17])
    SB_DFF i152_153 (.Q(ram_s_5_6), .C(CLK_3P3_MHZ_c), .D(n2982));   // src/ram.vhd(56[12:17])
    SB_DFF i149_150 (.Q(ram_s_5_5), .C(CLK_3P3_MHZ_c), .D(n2981));   // src/ram.vhd(56[12:17])
    SB_DFF i146_147 (.Q(ram_s_5_4), .C(CLK_3P3_MHZ_c), .D(n2980));   // src/ram.vhd(56[12:17])
    SB_DFF i143_144 (.Q(ram_s_5_3), .C(CLK_3P3_MHZ_c), .D(n2979));   // src/ram.vhd(56[12:17])
    SB_DFF i140_141 (.Q(ram_s_5_2), .C(CLK_3P3_MHZ_c), .D(n2978));   // src/ram.vhd(56[12:17])
    SB_DFF i137_138 (.Q(ram_s_5_1), .C(CLK_3P3_MHZ_c), .D(n2977));   // src/ram.vhd(56[12:17])
    SB_DFF i134_135 (.Q(ram_s_5_0), .C(CLK_3P3_MHZ_c), .D(n2976));   // src/ram.vhd(56[12:17])
    SB_DFF i131_132 (.Q(ram_s_4_7), .C(CLK_3P3_MHZ_c), .D(n2975));   // src/ram.vhd(56[12:17])
    SB_DFF i128_129 (.Q(ram_s_4_6), .C(CLK_3P3_MHZ_c), .D(n2974));   // src/ram.vhd(56[12:17])
    SB_DFF i125_126 (.Q(ram_s_4_5), .C(CLK_3P3_MHZ_c), .D(n2973));   // src/ram.vhd(56[12:17])
    SB_DFF i122_123 (.Q(ram_s_4_4), .C(CLK_3P3_MHZ_c), .D(n2972));   // src/ram.vhd(56[12:17])
    SB_DFF i119_120 (.Q(ram_s_4_3), .C(CLK_3P3_MHZ_c), .D(n2971));   // src/ram.vhd(56[12:17])
    SB_DFF i116_117 (.Q(ram_s_4_2), .C(CLK_3P3_MHZ_c), .D(n2970));   // src/ram.vhd(56[12:17])
    SB_DFF i113_114 (.Q(ram_s_4_1), .C(CLK_3P3_MHZ_c), .D(n2969));   // src/ram.vhd(56[12:17])
    SB_DFF i110_111 (.Q(ram_s_4_0), .C(CLK_3P3_MHZ_c), .D(n2968));   // src/ram.vhd(56[12:17])
    SB_DFF i107_108 (.Q(ram_s_3_7), .C(CLK_3P3_MHZ_c), .D(n2967));   // src/ram.vhd(56[12:17])
    SB_DFF i104_105 (.Q(ram_s_3_6), .C(CLK_3P3_MHZ_c), .D(n2966));   // src/ram.vhd(56[12:17])
    SB_DFF i101_102 (.Q(ram_s_3_5), .C(CLK_3P3_MHZ_c), .D(n2965));   // src/ram.vhd(56[12:17])
    SB_DFF i98_99 (.Q(ram_s_3_4), .C(CLK_3P3_MHZ_c), .D(n2964));   // src/ram.vhd(56[12:17])
    SB_DFF i95_96 (.Q(ram_s_3_3), .C(CLK_3P3_MHZ_c), .D(n2963));   // src/ram.vhd(56[12:17])
    SB_DFF i92_93 (.Q(ram_s_3_2), .C(CLK_3P3_MHZ_c), .D(n2962));   // src/ram.vhd(56[12:17])
    SB_DFF i89_90 (.Q(ram_s_3_1), .C(CLK_3P3_MHZ_c), .D(n2961));   // src/ram.vhd(56[12:17])
    SB_DFF i86_87 (.Q(ram_s_3_0), .C(CLK_3P3_MHZ_c), .D(n2960));   // src/ram.vhd(56[12:17])
    SB_DFF i83_84 (.Q(ram_s_2_7), .C(CLK_3P3_MHZ_c), .D(n2959));   // src/ram.vhd(56[12:17])
    SB_DFF i80_81 (.Q(ram_s_2_6), .C(CLK_3P3_MHZ_c), .D(n2958));   // src/ram.vhd(56[12:17])
    SB_DFF i77_78 (.Q(ram_s_2_5), .C(CLK_3P3_MHZ_c), .D(n2957));   // src/ram.vhd(56[12:17])
    SB_DFF i74_75 (.Q(ram_s_2_4), .C(CLK_3P3_MHZ_c), .D(n2956));   // src/ram.vhd(56[12:17])
    SB_DFF i71_72 (.Q(ram_s_2_3), .C(CLK_3P3_MHZ_c), .D(n2955));   // src/ram.vhd(56[12:17])
    SB_DFF i68_69 (.Q(ram_s_2_2), .C(CLK_3P3_MHZ_c), .D(n2954));   // src/ram.vhd(56[12:17])
    SB_DFF i65_66 (.Q(ram_s_2_1), .C(CLK_3P3_MHZ_c), .D(n2953));   // src/ram.vhd(56[12:17])
    SB_DFF i62_63 (.Q(ram_s_2_0), .C(CLK_3P3_MHZ_c), .D(n2952));   // src/ram.vhd(56[12:17])
    SB_DFF i59_60 (.Q(ram_s_1_7), .C(CLK_3P3_MHZ_c), .D(n2951));   // src/ram.vhd(56[12:17])
    SB_DFF i56_57 (.Q(ram_s_1_6), .C(CLK_3P3_MHZ_c), .D(n2950));   // src/ram.vhd(56[12:17])
    SB_DFF i53_54 (.Q(ram_s_1_5), .C(CLK_3P3_MHZ_c), .D(n2949));   // src/ram.vhd(56[12:17])
    SB_DFF i50_51 (.Q(ram_s_1_4), .C(CLK_3P3_MHZ_c), .D(n2948));   // src/ram.vhd(56[12:17])
    SB_DFF i47_48 (.Q(ram_s_1_3), .C(CLK_3P3_MHZ_c), .D(n2947));   // src/ram.vhd(56[12:17])
    SB_DFF i44_45 (.Q(ram_s_1_2), .C(CLK_3P3_MHZ_c), .D(n2946));   // src/ram.vhd(56[12:17])
    SB_DFF i41_42 (.Q(ram_s_1_1), .C(CLK_3P3_MHZ_c), .D(n2945));   // src/ram.vhd(56[12:17])
    SB_DFF i38_39 (.Q(ram_s_1_0), .C(CLK_3P3_MHZ_c), .D(n2944));   // src/ram.vhd(56[12:17])
    SB_DFF i35_36 (.Q(ram_s_0_7), .C(CLK_3P3_MHZ_c), .D(n2943));   // src/ram.vhd(56[12:17])
    SB_DFF i32_33 (.Q(ram_s_0_6), .C(CLK_3P3_MHZ_c), .D(n2942));   // src/ram.vhd(56[12:17])
    SB_DFF i29_30 (.Q(ram_s_0_5), .C(CLK_3P3_MHZ_c), .D(n2941));   // src/ram.vhd(56[12:17])
    SB_DFF i26_27 (.Q(ram_s_0_4), .C(CLK_3P3_MHZ_c), .D(n2940));   // src/ram.vhd(56[12:17])
    SB_DFF i23_24 (.Q(ram_s_0_3), .C(CLK_3P3_MHZ_c), .D(n2939));   // src/ram.vhd(56[12:17])
    SB_DFF i20_21 (.Q(ram_s_0_2), .C(CLK_3P3_MHZ_c), .D(n2938));   // src/ram.vhd(56[12:17])
    SB_DFF i17_18 (.Q(ram_s_0_1), .C(CLK_3P3_MHZ_c), .D(n2937));   // src/ram.vhd(56[12:17])
    SB_DFF i14_15 (.Q(ram_s_0_0), .C(CLK_3P3_MHZ_c), .D(n2936));   // src/ram.vhd(56[12:17])
    SB_LUT4 instruction_8__bdd_4_lut_10372 (.I0(\instruction[8] ), .I1(ram_s_6_5), 
            .I2(ram_s_7_5), .I3(\instruction[9] ), .O(n11471));
    defparam instruction_8__bdd_4_lut_10372.LUT_INIT = 16'he4aa;
    SB_LUT4 n11471_bdd_4_lut (.I0(n11471), .I1(ram_s_5_5), .I2(ram_s_4_5), 
            .I3(\instruction[9] ), .O(n11474));
    defparam n11471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10357 (.I0(\instruction[8] ), .I1(ram_s_22_3), 
            .I2(ram_s_23_3), .I3(\instruction[9] ), .O(n11435));
    defparam instruction_8__bdd_4_lut_10357.LUT_INIT = 16'he4aa;
    SB_LUT4 n11435_bdd_4_lut (.I0(n11435), .I1(ram_s_21_3), .I2(ram_s_20_3), 
            .I3(\instruction[9] ), .O(n11438));
    defparam n11435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_9__bdd_4_lut_11813 (.I0(\instruction[9] ), .I1(n8826), 
            .I2(n8827), .I3(\instruction[10] ), .O(n11345));
    defparam instruction_9__bdd_4_lut_11813.LUT_INIT = 16'he4aa;
    SB_LUT4 n11345_bdd_4_lut (.I0(n11345), .I1(n8809), .I2(n8808), .I3(\instruction[10] ), 
            .O(n11348));
    defparam n11345_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_9__bdd_4_lut_10253 (.I0(\instruction[9] ), .I1(n9657), 
            .I2(n9658), .I3(\instruction[10] ), .O(n11339));
    defparam instruction_9__bdd_4_lut_10253.LUT_INIT = 16'he4aa;
    SB_LUT4 n11339_bdd_4_lut (.I0(n11339), .I1(n9280), .I2(n9279), .I3(\instruction[10] ), 
            .O(n11342));
    defparam n11339_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_11__bdd_4_lut_10785 (.I0(\instruction[11] ), .I1(n11264), 
            .I2(n8806), .I3(\sx_addr[4] ), .O(n11315));
    defparam instruction_11__bdd_4_lut_10785.LUT_INIT = 16'he4aa;
    SB_LUT4 n11315_bdd_4_lut (.I0(n11315), .I1(n8800), .I2(n11234), .I3(\sx_addr[4] ), 
            .O(\register_vector[9] ));
    defparam n11315_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10328 (.I0(\instruction[8] ), .I1(ram_s_10_6), 
            .I2(ram_s_11_6), .I3(\instruction[9] ), .O(n11303));
    defparam instruction_8__bdd_4_lut_10328.LUT_INIT = 16'he4aa;
    SB_LUT4 n11303_bdd_4_lut (.I0(n11303), .I1(ram_s_9_6), .I2(ram_s_8_6), 
            .I3(\instruction[9] ), .O(n11306));
    defparam n11303_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10219 (.I0(\instruction[8] ), .I1(ram_s_30_6), 
            .I2(ram_s_31_6), .I3(\instruction[9] ), .O(n11273));
    defparam instruction_8__bdd_4_lut_10219.LUT_INIT = 16'he4aa;
    SB_LUT4 n11273_bdd_4_lut (.I0(n11273), .I1(ram_s_29_6), .I2(ram_s_28_6), 
            .I3(\instruction[9] ), .O(n11276));
    defparam n11273_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_9__bdd_4_lut_10248 (.I0(\instruction[9] ), .I1(n11073), 
            .I2(n11074), .I3(\instruction[10] ), .O(n11261));
    defparam instruction_9__bdd_4_lut_10248.LUT_INIT = 16'he4aa;
    SB_LUT4 n11261_bdd_4_lut (.I0(n11261), .I1(n11065), .I2(n11064), .I3(\instruction[10] ), 
            .O(n11264));
    defparam n11261_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2944_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_31_7), .O(n3192));   // src/ram.vhd(68[19:45])
    defparam i2944_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2943_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_31_6), .O(n3191));   // src/ram.vhd(68[19:45])
    defparam i2943_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2942_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_31_5), .O(n3190));   // src/ram.vhd(68[19:45])
    defparam i2942_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2941_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_31_4), .O(n3189));   // src/ram.vhd(68[19:45])
    defparam i2941_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2940_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_31_3), .O(n3188));   // src/ram.vhd(68[19:45])
    defparam i2940_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2939_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_31_2), .O(n3187));   // src/ram.vhd(68[19:45])
    defparam i2939_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2938_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_31_1), .O(n3186));   // src/ram.vhd(68[19:45])
    defparam i2938_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2937_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_31_0), .O(n3185));   // src/ram.vhd(68[19:45])
    defparam i2937_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i26_2_lut_3_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n26));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i26_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i27_2_lut_3_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n27));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i27_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i2936_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_30_7), .O(n3184));   // src/ram.vhd(68[19:45])
    defparam i2936_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2935_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_30_6), .O(n3183));   // src/ram.vhd(68[19:45])
    defparam i2935_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2934_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_30_5), .O(n3182));   // src/ram.vhd(68[19:45])
    defparam i2934_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2933_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_30_4), .O(n3181));   // src/ram.vhd(68[19:45])
    defparam i2933_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2932_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_30_3), .O(n3180));   // src/ram.vhd(68[19:45])
    defparam i2932_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2931_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_30_2), .O(n3179));   // src/ram.vhd(68[19:45])
    defparam i2931_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2930_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_30_1), .O(n3178));   // src/ram.vhd(68[19:45])
    defparam i2930_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2929_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_30_0), .O(n3177));   // src/ram.vhd(68[19:45])
    defparam i2929_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i24_2_lut_3_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n24));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i24_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i25_2_lut_3_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n25));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i25_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i2928_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_29_7), .O(n3176));   // src/ram.vhd(68[19:45])
    defparam i2928_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2926_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_29_6), .O(n3174));   // src/ram.vhd(68[19:45])
    defparam i2926_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2925_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_29_5), .O(n3173));   // src/ram.vhd(68[19:45])
    defparam i2925_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2924_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_29_4), .O(n3172));   // src/ram.vhd(68[19:45])
    defparam i2924_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2923_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_29_3), .O(n3171));   // src/ram.vhd(68[19:45])
    defparam i2923_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2922_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_29_2), .O(n3170));   // src/ram.vhd(68[19:45])
    defparam i2922_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2921_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_29_1), .O(n3169));   // src/ram.vhd(68[19:45])
    defparam i2921_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2920_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_29_0), .O(n3168));   // src/ram.vhd(68[19:45])
    defparam i2920_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i22_2_lut_3_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n22));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i22_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i23_2_lut_3_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n23));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i23_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i415630_i1_3_lut (.I0(n11918), .I1(n11906), .I2(\sx_addr[4] ), 
            .I3(wea[0]), .O(\register_vector[8] ));
    defparam i415630_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7762_3_lut (.I0(n13040), .I1(n12980), .I2(\instruction[10] ), 
            .I3(wea[0]), .O(n8821));
    defparam i7762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7763_3_lut (.I0(n11348), .I1(n8821), .I2(\instruction[11] ), 
            .I3(wea[0]), .O(n8822));
    defparam i7763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i420454_i1_3_lut (.I0(n8822), .I1(n11552), .I2(\sx_addr[4] ), 
            .I3(wea[0]), .O(\register_vector[10] ));
    defparam i420454_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i425278_i1_3_lut (.I0(n14786), .I1(n13748), .I2(\sx_addr[4] ), 
            .I3(wea[0]), .O(\sx[4] ));
    defparam i425278_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i427690_i1_3_lut (.I0(n11654), .I1(n12200), .I2(\sx_addr[4] ), 
            .I3(wea[0]), .O(\sx[5] ));
    defparam i427690_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4300102_i1_3_lut (.I0(n14378), .I1(n12374), .I2(\sx_addr[4] ), 
            .I3(wea[0]), .O(\sx[6] ));
    defparam i4300102_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4324114_i1_3_lut (.I0(n12206), .I1(n12548), .I2(\sx_addr[4] ), 
            .I3(wea[0]), .O(\sx[7] ));
    defparam i4324114_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2919_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_28_7), .O(n3167));   // src/ram.vhd(68[19:45])
    defparam i2919_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2918_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_28_6), .O(n3166));   // src/ram.vhd(68[19:45])
    defparam i2918_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2917_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_28_5), .O(n3165));   // src/ram.vhd(68[19:45])
    defparam i2917_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2916_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_28_4), .O(n3164));   // src/ram.vhd(68[19:45])
    defparam i2916_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2915_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_28_3), .O(n3163));   // src/ram.vhd(68[19:45])
    defparam i2915_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2914_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_28_2), .O(n3162));   // src/ram.vhd(68[19:45])
    defparam i2914_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2913_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_28_1), .O(n3161));   // src/ram.vhd(68[19:45])
    defparam i2913_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2912_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_28_0), .O(n3160));   // src/ram.vhd(68[19:45])
    defparam i2912_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i20_2_lut_3_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n20));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i20_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i21_2_lut_3_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[11] ), .I3(\instruction[10] ), .O(n21));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i21_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i2911_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_27_7), .O(n3159));   // src/ram.vhd(68[19:45])
    defparam i2911_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2910_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_27_6), .O(n3158));   // src/ram.vhd(68[19:45])
    defparam i2910_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2909_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_27_5), .O(n3157));   // src/ram.vhd(68[19:45])
    defparam i2909_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2908_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_27_4), .O(n3156));   // src/ram.vhd(68[19:45])
    defparam i2908_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2907_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_27_3), .O(n3155));   // src/ram.vhd(68[19:45])
    defparam i2907_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2906_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_27_2), .O(n3154));   // src/ram.vhd(68[19:45])
    defparam i2906_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2905_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_27_1), .O(n3153));   // src/ram.vhd(68[19:45])
    defparam i2905_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2904_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_27_0), .O(n3152));   // src/ram.vhd(68[19:45])
    defparam i2904_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2903_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_26_7), .O(n3151));   // src/ram.vhd(68[19:45])
    defparam i2903_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2902_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_26_6), .O(n3150));   // src/ram.vhd(68[19:45])
    defparam i2902_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2901_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_26_5), .O(n3149));   // src/ram.vhd(68[19:45])
    defparam i2901_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2900_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_26_4), .O(n3148));   // src/ram.vhd(68[19:45])
    defparam i2900_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2899_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_26_3), .O(n3147));   // src/ram.vhd(68[19:45])
    defparam i2899_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2898_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_26_2), .O(n3146));   // src/ram.vhd(68[19:45])
    defparam i2898_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2897_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_26_1), .O(n3145));   // src/ram.vhd(68[19:45])
    defparam i2897_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2896_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_26_0), .O(n3144));   // src/ram.vhd(68[19:45])
    defparam i2896_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2895_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_25_7), .O(n3143));   // src/ram.vhd(68[19:45])
    defparam i2895_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2894_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_25_6), .O(n3142));   // src/ram.vhd(68[19:45])
    defparam i2894_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2893_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_25_5), .O(n3141));   // src/ram.vhd(68[19:45])
    defparam i2893_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i29_2_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n29));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i29_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i28_2_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n28));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i28_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i2892_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_25_4), .O(n3140));   // src/ram.vhd(68[19:45])
    defparam i2892_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2891_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_25_3), .O(n3139));   // src/ram.vhd(68[19:45])
    defparam i2891_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2890_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_25_2), .O(n3138));   // src/ram.vhd(68[19:45])
    defparam i2890_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2889_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_25_1), .O(n3137));   // src/ram.vhd(68[19:45])
    defparam i2889_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2888_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_25_0), .O(n3136));   // src/ram.vhd(68[19:45])
    defparam i2888_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2887_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_24_7), .O(n3135));   // src/ram.vhd(68[19:45])
    defparam i2887_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2886_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_24_6), .O(n3134));   // src/ram.vhd(68[19:45])
    defparam i2886_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2885_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_24_5), .O(n3133));   // src/ram.vhd(68[19:45])
    defparam i2885_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2884_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_24_4), .O(n3132));   // src/ram.vhd(68[19:45])
    defparam i2884_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2883_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_24_3), .O(n3131));   // src/ram.vhd(68[19:45])
    defparam i2883_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2882_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_24_2), .O(n3130));   // src/ram.vhd(68[19:45])
    defparam i2882_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2881_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_24_1), .O(n3129));   // src/ram.vhd(68[19:45])
    defparam i2881_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2880_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_24_0), .O(n3128));   // src/ram.vhd(68[19:45])
    defparam i2880_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2879_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_23_7), .O(n3127));   // src/ram.vhd(68[19:45])
    defparam i2879_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2878_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_23_6), .O(n3126));   // src/ram.vhd(68[19:45])
    defparam i2878_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2877_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_23_5), .O(n3125));   // src/ram.vhd(68[19:45])
    defparam i2877_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2876_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_23_4), .O(n3124));   // src/ram.vhd(68[19:45])
    defparam i2876_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2875_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_23_3), .O(n3123));   // src/ram.vhd(68[19:45])
    defparam i2875_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2874_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_23_2), .O(n3122));   // src/ram.vhd(68[19:45])
    defparam i2874_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2873_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_23_1), .O(n3121));   // src/ram.vhd(68[19:45])
    defparam i2873_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2872_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_23_0), .O(n3120));   // src/ram.vhd(68[19:45])
    defparam i2872_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i7_2_lut (.I0(register_enable), .I1(\instruction[8] ), 
            .I2(wea[0]), .I3(wea[0]), .O(n7));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i7_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2871_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_22_7), .O(n3119));   // src/ram.vhd(68[19:45])
    defparam i2871_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2870_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_22_6), .O(n3118));   // src/ram.vhd(68[19:45])
    defparam i2870_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2869_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_22_5), .O(n3117));   // src/ram.vhd(68[19:45])
    defparam i2869_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2868_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_22_4), .O(n3116));   // src/ram.vhd(68[19:45])
    defparam i2868_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2867_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_22_3), .O(n3115));   // src/ram.vhd(68[19:45])
    defparam i2867_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2866_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_22_2), .O(n3114));   // src/ram.vhd(68[19:45])
    defparam i2866_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2865_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_22_1), .O(n3113));   // src/ram.vhd(68[19:45])
    defparam i2865_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2864_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_22_0), .O(n3112));   // src/ram.vhd(68[19:45])
    defparam i2864_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2863_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_21_7), .O(n3111));   // src/ram.vhd(68[19:45])
    defparam i2863_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2862_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_21_6), .O(n3110));   // src/ram.vhd(68[19:45])
    defparam i2862_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2861_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_21_5), .O(n3109));   // src/ram.vhd(68[19:45])
    defparam i2861_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2860_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_21_4), .O(n3108));   // src/ram.vhd(68[19:45])
    defparam i2860_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2859_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_21_3), .O(n3107));   // src/ram.vhd(68[19:45])
    defparam i2859_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2858_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_21_2), .O(n3106));   // src/ram.vhd(68[19:45])
    defparam i2858_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2857_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_21_1), .O(n3105));   // src/ram.vhd(68[19:45])
    defparam i2857_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2856_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_21_0), .O(n3104));   // src/ram.vhd(68[19:45])
    defparam i2856_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2855_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_20_7), .O(n3103));   // src/ram.vhd(68[19:45])
    defparam i2855_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2854_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_20_6), .O(n3102));   // src/ram.vhd(68[19:45])
    defparam i2854_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2853_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_20_5), .O(n3101));   // src/ram.vhd(68[19:45])
    defparam i2853_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2852_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_20_4), .O(n3100));   // src/ram.vhd(68[19:45])
    defparam i2852_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2851_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_20_3), .O(n3099));   // src/ram.vhd(68[19:45])
    defparam i2851_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2850_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_20_2), .O(n3098));   // src/ram.vhd(68[19:45])
    defparam i2850_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2849_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_20_1), .O(n3097));   // src/ram.vhd(68[19:45])
    defparam i2849_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2848_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_20_0), .O(n3096));   // src/ram.vhd(68[19:45])
    defparam i2848_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2847_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_19_7), .O(n3095));   // src/ram.vhd(68[19:45])
    defparam i2847_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2846_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_19_6), .O(n3094));   // src/ram.vhd(68[19:45])
    defparam i2846_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2845_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_19_5), .O(n3093));   // src/ram.vhd(68[19:45])
    defparam i2845_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2844_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_19_4), .O(n3092));   // src/ram.vhd(68[19:45])
    defparam i2844_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2843_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_19_3), .O(n3091));   // src/ram.vhd(68[19:45])
    defparam i2843_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2842_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_19_2), .O(n3090));   // src/ram.vhd(68[19:45])
    defparam i2842_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2841_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_19_1), .O(n3089));   // src/ram.vhd(68[19:45])
    defparam i2841_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2840_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_19_0), .O(n3088));   // src/ram.vhd(68[19:45])
    defparam i2840_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2839_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_18_7), .O(n3087));   // src/ram.vhd(68[19:45])
    defparam i2839_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2838_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_18_6), .O(n3086));   // src/ram.vhd(68[19:45])
    defparam i2838_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2837_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_18_5), .O(n3085));   // src/ram.vhd(68[19:45])
    defparam i2837_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2836_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_18_4), .O(n3084));   // src/ram.vhd(68[19:45])
    defparam i2836_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2835_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_18_3), .O(n3083));   // src/ram.vhd(68[19:45])
    defparam i2835_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2834_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_18_2), .O(n3082));   // src/ram.vhd(68[19:45])
    defparam i2834_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2833_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_18_1), .O(n3081));   // src/ram.vhd(68[19:45])
    defparam i2833_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2832_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_18_0), .O(n3080));   // src/ram.vhd(68[19:45])
    defparam i2832_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2831_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_17_7), .O(n3079));   // src/ram.vhd(68[19:45])
    defparam i2831_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2830_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_17_6), .O(n3078));   // src/ram.vhd(68[19:45])
    defparam i2830_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2829_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_17_5), .O(n3077));   // src/ram.vhd(68[19:45])
    defparam i2829_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2828_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_17_4), .O(n3076));   // src/ram.vhd(68[19:45])
    defparam i2828_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2827_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_17_3), .O(n3075));   // src/ram.vhd(68[19:45])
    defparam i2827_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2826_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_17_2), .O(n3074));   // src/ram.vhd(68[19:45])
    defparam i2826_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2825_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_17_1), .O(n3073));   // src/ram.vhd(68[19:45])
    defparam i2825_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2824_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_17_0), .O(n3072));   // src/ram.vhd(68[19:45])
    defparam i2824_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i31_2_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n31));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i31_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i2823_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_16_7), .O(n3071));   // src/ram.vhd(68[19:45])
    defparam i2823_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2822_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_16_6), .O(n3070));   // src/ram.vhd(68[19:45])
    defparam i2822_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2821_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_16_5), .O(n3069));   // src/ram.vhd(68[19:45])
    defparam i2821_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2820_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_16_4), .O(n3068));   // src/ram.vhd(68[19:45])
    defparam i2820_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2819_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_16_3), .O(n3067));   // src/ram.vhd(68[19:45])
    defparam i2819_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2818_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_16_2), .O(n3066));   // src/ram.vhd(68[19:45])
    defparam i2818_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2817_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_16_1), .O(n3065));   // src/ram.vhd(68[19:45])
    defparam i2817_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2816_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_16_0), .O(n3064));   // src/ram.vhd(68[19:45])
    defparam i2816_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2815_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_15_7), .O(n3063));   // src/ram.vhd(68[19:45])
    defparam i2815_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2814_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_15_6), .O(n3062));   // src/ram.vhd(68[19:45])
    defparam i2814_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2813_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_15_5), .O(n3061));   // src/ram.vhd(68[19:45])
    defparam i2813_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2812_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_15_4), .O(n3060));   // src/ram.vhd(68[19:45])
    defparam i2812_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2811_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_15_3), .O(n3059));   // src/ram.vhd(68[19:45])
    defparam i2811_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2810_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_15_2), .O(n3058));   // src/ram.vhd(68[19:45])
    defparam i2810_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2809_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_15_1), .O(n3057));   // src/ram.vhd(68[19:45])
    defparam i2809_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2808_3_lut_4_lut (.I0(n34), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_15_0), .O(n3056));   // src/ram.vhd(68[19:45])
    defparam i2808_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2807_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_14_7), .O(n3055));   // src/ram.vhd(68[19:45])
    defparam i2807_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2806_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_14_6), .O(n3054));   // src/ram.vhd(68[19:45])
    defparam i2806_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2805_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_14_5), .O(n3053));   // src/ram.vhd(68[19:45])
    defparam i2805_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2804_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_14_4), .O(n3052));   // src/ram.vhd(68[19:45])
    defparam i2804_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2803_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_14_3), .O(n3051));   // src/ram.vhd(68[19:45])
    defparam i2803_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2802_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_14_2), .O(n3050));   // src/ram.vhd(68[19:45])
    defparam i2802_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2801_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_14_1), .O(n3049));   // src/ram.vhd(68[19:45])
    defparam i2801_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2800_3_lut_4_lut (.I0(n32), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_14_0), .O(n3048));   // src/ram.vhd(68[19:45])
    defparam i2800_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2799_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_13_7), .O(n3047));   // src/ram.vhd(68[19:45])
    defparam i2799_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2798_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_13_6), .O(n3046));   // src/ram.vhd(68[19:45])
    defparam i2798_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2797_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_13_5), .O(n3045));   // src/ram.vhd(68[19:45])
    defparam i2797_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2796_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_13_4), .O(n3044));   // src/ram.vhd(68[19:45])
    defparam i2796_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2795_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_13_3), .O(n3043));   // src/ram.vhd(68[19:45])
    defparam i2795_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2794_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_13_2), .O(n3042));   // src/ram.vhd(68[19:45])
    defparam i2794_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2793_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_13_1), .O(n3041));   // src/ram.vhd(68[19:45])
    defparam i2793_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2792_3_lut_4_lut (.I0(n30), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_13_0), .O(n3040));   // src/ram.vhd(68[19:45])
    defparam i2792_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2791_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_12_7), .O(n3039));   // src/ram.vhd(68[19:45])
    defparam i2791_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2790_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_12_6), .O(n3038));   // src/ram.vhd(68[19:45])
    defparam i2790_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2789_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_12_5), .O(n3037));   // src/ram.vhd(68[19:45])
    defparam i2789_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2788_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_12_4), .O(n3036));   // src/ram.vhd(68[19:45])
    defparam i2788_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2787_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_12_3), .O(n3035));   // src/ram.vhd(68[19:45])
    defparam i2787_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2786_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_12_2), .O(n3034));   // src/ram.vhd(68[19:45])
    defparam i2786_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2785_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_12_1), .O(n3033));   // src/ram.vhd(68[19:45])
    defparam i2785_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2784_3_lut_4_lut (.I0(n28), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_12_0), .O(n3032));   // src/ram.vhd(68[19:45])
    defparam i2784_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2783_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_11_7), .O(n3031));   // src/ram.vhd(68[19:45])
    defparam i2783_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2782_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_11_6), .O(n3030));   // src/ram.vhd(68[19:45])
    defparam i2782_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2781_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_11_5), .O(n3029));   // src/ram.vhd(68[19:45])
    defparam i2781_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2780_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_11_4), .O(n3028));   // src/ram.vhd(68[19:45])
    defparam i2780_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2779_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_11_3), .O(n3027));   // src/ram.vhd(68[19:45])
    defparam i2779_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2778_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_11_2), .O(n3026));   // src/ram.vhd(68[19:45])
    defparam i2778_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2777_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_11_1), .O(n3025));   // src/ram.vhd(68[19:45])
    defparam i2777_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2776_3_lut_4_lut (.I0(n26), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_11_0), .O(n3024));   // src/ram.vhd(68[19:45])
    defparam i2776_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2775_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_10_7), .O(n3023));   // src/ram.vhd(68[19:45])
    defparam i2775_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2774_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_10_6), .O(n3022));   // src/ram.vhd(68[19:45])
    defparam i2774_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2773_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_10_5), .O(n3021));   // src/ram.vhd(68[19:45])
    defparam i2773_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2772_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_10_4), .O(n3020));   // src/ram.vhd(68[19:45])
    defparam i2772_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2771_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_10_3), .O(n3019));   // src/ram.vhd(68[19:45])
    defparam i2771_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2770_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_10_2), .O(n3018));   // src/ram.vhd(68[19:45])
    defparam i2770_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2769_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_10_1), .O(n3017));   // src/ram.vhd(68[19:45])
    defparam i2769_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2768_3_lut_4_lut (.I0(n24), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_10_0), .O(n3016));   // src/ram.vhd(68[19:45])
    defparam i2768_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2767_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_9_7), .O(n3015));   // src/ram.vhd(68[19:45])
    defparam i2767_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2766_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_9_6), .O(n3014));   // src/ram.vhd(68[19:45])
    defparam i2766_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2765_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_9_5), .O(n3013));   // src/ram.vhd(68[19:45])
    defparam i2765_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2764_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_9_4), .O(n3012));   // src/ram.vhd(68[19:45])
    defparam i2764_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2763_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_9_3), .O(n3011));   // src/ram.vhd(68[19:45])
    defparam i2763_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2762_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_9_2), .O(n3010));   // src/ram.vhd(68[19:45])
    defparam i2762_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2761_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_9_1), .O(n3009));   // src/ram.vhd(68[19:45])
    defparam i2761_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2760_3_lut_4_lut (.I0(n22), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_9_0), .O(n3008));   // src/ram.vhd(68[19:45])
    defparam i2760_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2759_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_8_7), .O(n3007));   // src/ram.vhd(68[19:45])
    defparam i2759_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2758_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_8_6), .O(n3006));   // src/ram.vhd(68[19:45])
    defparam i2758_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2757_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_8_5), .O(n3005));   // src/ram.vhd(68[19:45])
    defparam i2757_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2756_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_8_4), .O(n3004));   // src/ram.vhd(68[19:45])
    defparam i2756_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2755_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_8_3), .O(n3003));   // src/ram.vhd(68[19:45])
    defparam i2755_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2754_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_8_2), .O(n3002));   // src/ram.vhd(68[19:45])
    defparam i2754_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2753_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_8_1), .O(n3001));   // src/ram.vhd(68[19:45])
    defparam i2753_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2752_3_lut_4_lut (.I0(n20), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_8_0), .O(n3000));   // src/ram.vhd(68[19:45])
    defparam i2752_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2751_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_7_7), .O(n2999));   // src/ram.vhd(68[19:45])
    defparam i2751_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2750_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_7_6), .O(n2998));   // src/ram.vhd(68[19:45])
    defparam i2750_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2749_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_7_5), .O(n2997));   // src/ram.vhd(68[19:45])
    defparam i2749_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2748_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_7_4), .O(n2996));   // src/ram.vhd(68[19:45])
    defparam i2748_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2747_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_7_3), .O(n2995));   // src/ram.vhd(68[19:45])
    defparam i2747_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2746_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_7_2), .O(n2994));   // src/ram.vhd(68[19:45])
    defparam i2746_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2745_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_7_1), .O(n2993));   // src/ram.vhd(68[19:45])
    defparam i2745_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2744_3_lut_4_lut (.I0(n35), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_7_0), .O(n2992));   // src/ram.vhd(68[19:45])
    defparam i2744_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2743_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_6_7), .O(n2991));   // src/ram.vhd(68[19:45])
    defparam i2743_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2742_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_6_6), .O(n2990));   // src/ram.vhd(68[19:45])
    defparam i2742_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2741_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_6_5), .O(n2989));   // src/ram.vhd(68[19:45])
    defparam i2741_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2740_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_6_4), .O(n2988));   // src/ram.vhd(68[19:45])
    defparam i2740_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2739_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_6_3), .O(n2987));   // src/ram.vhd(68[19:45])
    defparam i2739_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2738_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_6_2), .O(n2986));   // src/ram.vhd(68[19:45])
    defparam i2738_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2737_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_6_1), .O(n2985));   // src/ram.vhd(68[19:45])
    defparam i2737_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2736_3_lut_4_lut (.I0(n33), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_6_0), .O(n2984));   // src/ram.vhd(68[19:45])
    defparam i2736_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2735_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_5_7), .O(n2983));   // src/ram.vhd(68[19:45])
    defparam i2735_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2734_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_5_6), .O(n2982));   // src/ram.vhd(68[19:45])
    defparam i2734_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2733_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_5_5), .O(n2981));   // src/ram.vhd(68[19:45])
    defparam i2733_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2732_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_5_4), .O(n2980));   // src/ram.vhd(68[19:45])
    defparam i2732_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2731_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_5_3), .O(n2979));   // src/ram.vhd(68[19:45])
    defparam i2731_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2730_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_5_2), .O(n2978));   // src/ram.vhd(68[19:45])
    defparam i2730_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2729_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_5_1), .O(n2977));   // src/ram.vhd(68[19:45])
    defparam i2729_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2728_3_lut_4_lut (.I0(n31), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_5_0), .O(n2976));   // src/ram.vhd(68[19:45])
    defparam i2728_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2727_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_4_7), .O(n2975));   // src/ram.vhd(68[19:45])
    defparam i2727_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2726_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_4_6), .O(n2974));   // src/ram.vhd(68[19:45])
    defparam i2726_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2725_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_4_5), .O(n2973));   // src/ram.vhd(68[19:45])
    defparam i2725_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2724_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_4_4), .O(n2972));   // src/ram.vhd(68[19:45])
    defparam i2724_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2723_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_4_3), .O(n2971));   // src/ram.vhd(68[19:45])
    defparam i2723_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2722_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_4_2), .O(n2970));   // src/ram.vhd(68[19:45])
    defparam i2722_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2721_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_4_1), .O(n2969));   // src/ram.vhd(68[19:45])
    defparam i2721_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2720_3_lut_4_lut (.I0(n29), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_4_0), .O(n2968));   // src/ram.vhd(68[19:45])
    defparam i2720_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2719_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_3_7), .O(n2967));   // src/ram.vhd(68[19:45])
    defparam i2719_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2718_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_3_6), .O(n2966));   // src/ram.vhd(68[19:45])
    defparam i2718_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2717_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_3_5), .O(n2965));   // src/ram.vhd(68[19:45])
    defparam i2717_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2716_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_3_4), .O(n2964));   // src/ram.vhd(68[19:45])
    defparam i2716_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2715_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_3_3), .O(n2963));   // src/ram.vhd(68[19:45])
    defparam i2715_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2714_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_3_2), .O(n2962));   // src/ram.vhd(68[19:45])
    defparam i2714_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2713_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_3_1), .O(n2961));   // src/ram.vhd(68[19:45])
    defparam i2713_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2712_3_lut_4_lut (.I0(n27), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_3_0), .O(n2960));   // src/ram.vhd(68[19:45])
    defparam i2712_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2711_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_2_7), .O(n2959));   // src/ram.vhd(68[19:45])
    defparam i2711_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2710_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_2_6), .O(n2958));   // src/ram.vhd(68[19:45])
    defparam i2710_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2709_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_2_5), .O(n2957));   // src/ram.vhd(68[19:45])
    defparam i2709_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2708_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_2_4), .O(n2956));   // src/ram.vhd(68[19:45])
    defparam i2708_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2707_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_2_3), .O(n2955));   // src/ram.vhd(68[19:45])
    defparam i2707_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2706_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_2_2), .O(n2954));   // src/ram.vhd(68[19:45])
    defparam i2706_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2705_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_2_1), .O(n2953));   // src/ram.vhd(68[19:45])
    defparam i2705_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2704_3_lut_4_lut (.I0(n25), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_2_0), .O(n2952));   // src/ram.vhd(68[19:45])
    defparam i2704_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2703_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_1_7), .O(n2951));   // src/ram.vhd(68[19:45])
    defparam i2703_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2702_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_1_6), .O(n2950));   // src/ram.vhd(68[19:45])
    defparam i2702_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2701_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_1_5), .O(n2949));   // src/ram.vhd(68[19:45])
    defparam i2701_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2700_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_1_4), .O(n2948));   // src/ram.vhd(68[19:45])
    defparam i2700_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2699_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_1_3), .O(n2947));   // src/ram.vhd(68[19:45])
    defparam i2699_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2698_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_1_2), .O(n2946));   // src/ram.vhd(68[19:45])
    defparam i2698_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2697_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_1_1), .O(n2945));   // src/ram.vhd(68[19:45])
    defparam i2697_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2696_3_lut_4_lut (.I0(n23), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_1_0), .O(n2944));   // src/ram.vhd(68[19:45])
    defparam i2696_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2695_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[7]), 
            .I3(ram_s_0_7), .O(n2943));   // src/ram.vhd(68[19:45])
    defparam i2695_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2694_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[6]), 
            .I3(ram_s_0_6), .O(n2942));   // src/ram.vhd(68[19:45])
    defparam i2694_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2693_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[5]), 
            .I3(ram_s_0_5), .O(n2941));   // src/ram.vhd(68[19:45])
    defparam i2693_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2692_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[4]), 
            .I3(ram_s_0_4), .O(n2940));   // src/ram.vhd(68[19:45])
    defparam i2692_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2691_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[3]), 
            .I3(ram_s_0_3), .O(n2939));   // src/ram.vhd(68[19:45])
    defparam i2691_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2690_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[2]), 
            .I3(ram_s_0_2), .O(n2938));   // src/ram.vhd(68[19:45])
    defparam i2690_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2689_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[1]), 
            .I3(ram_s_0_1), .O(n2937));   // src/ram.vhd(68[19:45])
    defparam i2689_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2688_3_lut_4_lut (.I0(n21), .I1(\sx_addr[4] ), .I2(alu_result[0]), 
            .I3(ram_s_0_0), .O(n2936));   // src/ram.vhd(68[19:45])
    defparam i2688_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i6_2_lut (.I0(register_enable), .I1(\instruction[8] ), 
            .I2(wea[0]), .I3(wea[0]), .O(n6));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 instruction_8__bdd_4_lut_11563 (.I0(\instruction[8] ), .I1(ram_s_18_5), 
            .I2(ram_s_19_5), .I3(\instruction[9] ), .O(n12815));
    defparam instruction_8__bdd_4_lut_11563.LUT_INIT = 16'he4aa;
    SB_LUT4 n12815_bdd_4_lut (.I0(n12815), .I1(ram_s_17_5), .I2(ram_s_16_5), 
            .I3(\instruction[9] ), .O(n10823));
    defparam n12815_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11473 (.I0(\instruction[8] ), .I1(ram_s_10_4), 
            .I2(ram_s_11_4), .I3(\instruction[9] ), .O(n12725));
    defparam instruction_8__bdd_4_lut_11473.LUT_INIT = 16'he4aa;
    SB_LUT4 n12725_bdd_4_lut (.I0(n12725), .I1(ram_s_9_4), .I2(ram_s_8_4), 
            .I3(\instruction[9] ), .O(n12728));
    defparam n12725_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10710 (.I0(\instruction[8] ), .I1(ram_s_6_0), 
            .I2(ram_s_7_0), .I3(\instruction[9] ), .O(n11879));
    defparam instruction_8__bdd_4_lut_10710.LUT_INIT = 16'he4aa;
    SB_LUT4 n11879_bdd_4_lut (.I0(n11879), .I1(ram_s_5_0), .I2(ram_s_4_0), 
            .I3(\instruction[9] ), .O(n11882));
    defparam n11879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_10506 (.I0(\instruction[10] ), .I1(n8858), 
            .I2(n8867), .I3(\instruction[11] ), .O(n11549));
    defparam instruction_10__bdd_4_lut_10506.LUT_INIT = 16'he4aa;
    SB_LUT4 n11549_bdd_4_lut (.I0(n11549), .I1(n8846), .I2(n8840), .I3(\instruction[11] ), 
            .O(n11552));
    defparam n11549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9966_3_lut (.I0(ram_s_0_1), .I1(ram_s_1_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11025));
    defparam i9966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9967_3_lut (.I0(ram_s_2_1), .I1(ram_s_3_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11026));
    defparam i9967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 instruction_8__bdd_4_lut_10695 (.I0(\instruction[8] ), .I1(ram_s_10_1), 
            .I2(ram_s_11_1), .I3(\instruction[9] ), .O(n11861));
    defparam instruction_8__bdd_4_lut_10695.LUT_INIT = 16'he4aa;
    SB_LUT4 n11861_bdd_4_lut (.I0(n11861), .I1(ram_s_9_1), .I2(ram_s_8_1), 
            .I3(\instruction[9] ), .O(n11864));
    defparam n11861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11398 (.I0(\instruction[8] ), .I1(ram_s_22_2), 
            .I2(ram_s_23_2), .I3(\instruction[9] ), .O(n12683));
    defparam instruction_8__bdd_4_lut_11398.LUT_INIT = 16'he4aa;
    SB_LUT4 n12683_bdd_4_lut (.I0(n12683), .I1(ram_s_21_2), .I2(ram_s_20_2), 
            .I3(\instruction[9] ), .O(n8846));
    defparam n12683_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10680 (.I0(\instruction[8] ), .I1(ram_s_10_0), 
            .I2(ram_s_11_0), .I3(\instruction[9] ), .O(n11843));
    defparam instruction_8__bdd_4_lut_10680.LUT_INIT = 16'he4aa;
    SB_LUT4 n11843_bdd_4_lut (.I0(n11843), .I1(ram_s_9_0), .I2(ram_s_8_0), 
            .I3(\instruction[9] ), .O(n11846));
    defparam n11843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9979_3_lut (.I0(ram_s_6_1), .I1(ram_s_7_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11038));
    defparam i9979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 instruction_8__bdd_4_lut_10581 (.I0(\instruction[8] ), .I1(ram_s_30_2), 
            .I2(ram_s_31_2), .I3(\instruction[9] ), .O(n11657));
    defparam instruction_8__bdd_4_lut_10581.LUT_INIT = 16'he4aa;
    SB_LUT4 i9978_3_lut (.I0(ram_s_4_1), .I1(ram_s_5_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11037));
    defparam i9978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 instruction_8__bdd_4_lut_10665 (.I0(\instruction[8] ), .I1(ram_s_14_1), 
            .I2(ram_s_15_1), .I3(\instruction[9] ), .O(n11831));
    defparam instruction_8__bdd_4_lut_10665.LUT_INIT = 16'he4aa;
    SB_LUT4 n11657_bdd_4_lut (.I0(n11657), .I1(ram_s_29_2), .I2(ram_s_28_2), 
            .I3(\instruction[9] ), .O(n8867));
    defparam n11657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11831_bdd_4_lut (.I0(n11831), .I1(ram_s_13_1), .I2(ram_s_12_1), 
            .I3(\instruction[9] ), .O(n11834));
    defparam n11831_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_10715 (.I0(\instruction[10] ), .I1(n10643), 
            .I2(n10733), .I3(\instruction[11] ), .O(n11651));
    defparam instruction_10__bdd_4_lut_10715.LUT_INIT = 16'he4aa;
    SB_LUT4 n11651_bdd_4_lut (.I0(n11651), .I1(n11474), .I2(n10466), .I3(\instruction[11] ), 
            .O(n11654));
    defparam n11651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10655 (.I0(\instruction[8] ), .I1(ram_s_14_0), 
            .I2(ram_s_15_0), .I3(\instruction[9] ), .O(n11825));
    defparam instruction_8__bdd_4_lut_10655.LUT_INIT = 16'he4aa;
    SB_LUT4 n11825_bdd_4_lut (.I0(n11825), .I1(ram_s_13_0), .I2(ram_s_12_0), 
            .I3(\instruction[9] ), .O(n11828));
    defparam n11825_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10511 (.I0(\instruction[8] ), .I1(ram_s_30_4), 
            .I2(ram_s_31_4), .I3(\instruction[9] ), .O(n11645));
    defparam instruction_8__bdd_4_lut_10511.LUT_INIT = 16'he4aa;
    SB_LUT4 n11645_bdd_4_lut (.I0(n11645), .I1(ram_s_29_4), .I2(ram_s_28_4), 
            .I3(\instruction[9] ), .O(n11648));
    defparam n11645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_12247 (.I0(\instruction[10] ), .I1(n10400), 
            .I2(n10421), .I3(\instruction[11] ), .O(n12545));
    defparam instruction_10__bdd_4_lut_12247.LUT_INIT = 16'he4aa;
    SB_LUT4 n12545_bdd_4_lut (.I0(n12545), .I1(n10355), .I2(n10310), .I3(\instruction[11] ), 
            .O(n12548));
    defparam n12545_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_11__bdd_4_lut (.I0(\instruction[11] ), .I1(n8994), 
            .I2(n8995), .I3(\sx_addr[4] ), .O(n11987));
    defparam instruction_11__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n11987_bdd_4_lut (.I0(n11987), .I1(n8818), .I2(n11342), .I3(\sx_addr[4] ), 
            .O(\register_vector[11] ));
    defparam n11987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_11105 (.I0(\instruction[10] ), .I1(n10235), 
            .I2(n10262), .I3(\instruction[11] ), .O(n12203));
    defparam instruction_10__bdd_4_lut_11105.LUT_INIT = 16'he4aa;
    SB_LUT4 n12203_bdd_4_lut (.I0(n12203), .I1(n11762), .I2(n10127), .I3(\instruction[11] ), 
            .O(n12206));
    defparam n12203_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_10965 (.I0(\instruction[10] ), .I1(n11948), 
            .I2(n8948), .I3(\instruction[11] ), .O(n12197));
    defparam instruction_10__bdd_4_lut_10965.LUT_INIT = 16'he4aa;
    SB_LUT4 n13217_bdd_4_lut (.I0(n13217), .I1(ram_s_5_6), .I2(ram_s_4_6), 
            .I3(\instruction[9] ), .O(n13220));
    defparam n13217_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11848 (.I0(\instruction[8] ), .I1(ram_s_6_6), 
            .I2(ram_s_7_6), .I3(\instruction[9] ), .O(n13217));
    defparam instruction_8__bdd_4_lut_11848.LUT_INIT = 16'he4aa;
    SB_LUT4 n13223_bdd_4_lut (.I0(n13223), .I1(n10033), .I2(n10032), .I3(\instruction[10] ), 
            .O(n8818));
    defparam n13223_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_9__bdd_4_lut (.I0(\instruction[9] ), .I1(n10290), 
            .I2(n10291), .I3(\instruction[10] ), .O(n13223));
    defparam instruction_9__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 instruction_8__bdd_4_lut_11363 (.I0(\instruction[8] ), .I1(ram_s_2_7), 
            .I2(ram_s_3_7), .I3(\instruction[9] ), .O(n12467));
    defparam instruction_8__bdd_4_lut_11363.LUT_INIT = 16'he4aa;
    SB_LUT4 n12467_bdd_4_lut (.I0(n12467), .I1(ram_s_1_7), .I2(ram_s_0_7), 
            .I3(\instruction[9] ), .O(n10127));
    defparam n12467_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11184 (.I0(\instruction[8] ), .I1(ram_s_26_1), 
            .I2(ram_s_27_1), .I3(\instruction[9] ), .O(n12431));
    defparam instruction_8__bdd_4_lut_11184.LUT_INIT = 16'he4aa;
    SB_LUT4 n12197_bdd_4_lut (.I0(n12197), .I1(n12152), .I2(n10823), .I3(\instruction[11] ), 
            .O(n12200));
    defparam n12197_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10650 (.I0(\instruction[8] ), .I1(ram_s_6_7), 
            .I2(ram_s_7_7), .I3(\instruction[9] ), .O(n11759));
    defparam instruction_8__bdd_4_lut_10650.LUT_INIT = 16'he4aa;
    SB_LUT4 n12431_bdd_4_lut (.I0(n12431), .I1(ram_s_25_1), .I2(ram_s_24_1), 
            .I3(\instruction[9] ), .O(n12434));
    defparam n12431_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11154 (.I0(\instruction[8] ), .I1(ram_s_2_5), 
            .I2(ram_s_3_5), .I3(\instruction[9] ), .O(n12389));
    defparam instruction_8__bdd_4_lut_11154.LUT_INIT = 16'he4aa;
    SB_LUT4 n12389_bdd_4_lut (.I0(n12389), .I1(ram_s_1_5), .I2(ram_s_0_5), 
            .I3(\instruction[9] ), .O(n10466));
    defparam n12389_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11100 (.I0(\instruction[8] ), .I1(ram_s_22_5), 
            .I2(ram_s_23_5), .I3(\instruction[9] ), .O(n12149));
    defparam instruction_8__bdd_4_lut_11100.LUT_INIT = 16'he4aa;
    SB_LUT4 n12149_bdd_4_lut (.I0(n12149), .I1(ram_s_21_5), .I2(ram_s_20_5), 
            .I3(\instruction[9] ), .O(n12152));
    defparam n12149_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_10880 (.I0(\instruction[8] ), .I1(ram_s_26_5), 
            .I2(ram_s_27_5), .I3(\instruction[9] ), .O(n11945));
    defparam instruction_8__bdd_4_lut_10880.LUT_INIT = 16'he4aa;
    SB_LUT4 n11945_bdd_4_lut (.I0(n11945), .I1(ram_s_25_5), .I2(ram_s_24_5), 
            .I3(\instruction[9] ), .O(n11948));
    defparam n11945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11759_bdd_4_lut (.I0(n11759), .I1(ram_s_5_7), .I2(ram_s_4_7), 
            .I3(\instruction[9] ), .O(n11762));
    defparam n11759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_11248 (.I0(\instruction[10] ), .I1(n12368), 
            .I2(n11276), .I3(\instruction[11] ), .O(n12371));
    defparam instruction_10__bdd_4_lut_11248.LUT_INIT = 16'he4aa;
    SB_LUT4 n12371_bdd_4_lut (.I0(n12371), .I1(n9653), .I2(n9560), .I3(\instruction[11] ), 
            .O(n12374));
    defparam n12371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13265_bdd_4_lut (.I0(n13265), .I1(ram_s_17_4), .I2(ram_s_16_4), 
            .I3(\instruction[9] ), .O(n13268));
    defparam n13265_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_11853 (.I0(\instruction[8] ), .I1(ram_s_18_4), 
            .I2(ram_s_19_4), .I3(\instruction[9] ), .O(n13265));
    defparam instruction_8__bdd_4_lut_11853.LUT_INIT = 16'he4aa;
    SB_LUT4 n13271_bdd_4_lut (.I0(n13271), .I1(ram_s_21_6), .I2(ram_s_20_6), 
            .I3(\instruction[9] ), .O(n9653));
    defparam n13271_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12048 (.I0(\instruction[8] ), .I1(ram_s_22_6), 
            .I2(ram_s_23_6), .I3(\instruction[9] ), .O(n13271));
    defparam instruction_8__bdd_4_lut_12048.LUT_INIT = 16'he4aa;
    SB_LUT4 n13505_bdd_4_lut (.I0(n13505), .I1(ram_s_25_7), .I2(ram_s_24_7), 
            .I3(\instruction[9] ), .O(n10400));
    defparam n13505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12063 (.I0(\instruction[8] ), .I1(ram_s_26_7), 
            .I2(ram_s_27_7), .I3(\instruction[9] ), .O(n13505));
    defparam instruction_8__bdd_4_lut_12063.LUT_INIT = 16'he4aa;
    SB_LUT4 n13523_bdd_4_lut (.I0(n13523), .I1(ram_s_25_4), .I2(ram_s_24_4), 
            .I3(\instruction[9] ), .O(n13526));
    defparam n13523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12098 (.I0(\instruction[8] ), .I1(ram_s_26_4), 
            .I2(ram_s_27_4), .I3(\instruction[9] ), .O(n13523));
    defparam instruction_8__bdd_4_lut_12098.LUT_INIT = 16'he4aa;
    SB_LUT4 n13565_bdd_4_lut (.I0(n13565), .I1(ram_s_29_1), .I2(ram_s_28_1), 
            .I3(\instruction[9] ), .O(n13568));
    defparam n13565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12227 (.I0(\instruction[8] ), .I1(ram_s_30_1), 
            .I2(ram_s_31_1), .I3(\instruction[9] ), .O(n13565));
    defparam instruction_8__bdd_4_lut_12227.LUT_INIT = 16'he4aa;
    SB_LUT4 n13721_bdd_4_lut (.I0(n13721), .I1(ram_s_17_3), .I2(ram_s_16_3), 
            .I3(\instruction[9] ), .O(n13724));
    defparam n13721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12242 (.I0(\instruction[8] ), .I1(ram_s_18_3), 
            .I2(ram_s_19_3), .I3(\instruction[9] ), .O(n13721));
    defparam instruction_8__bdd_4_lut_12242.LUT_INIT = 16'he4aa;
    SB_LUT4 n13739_bdd_4_lut (.I0(n13739), .I1(ram_s_25_3), .I2(ram_s_24_3), 
            .I3(\instruction[9] ), .O(n13742));
    defparam n13739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12252 (.I0(\instruction[8] ), .I1(ram_s_26_3), 
            .I2(ram_s_27_3), .I3(\instruction[9] ), .O(n13739));
    defparam instruction_8__bdd_4_lut_12252.LUT_INIT = 16'he4aa;
    SB_LUT4 n13745_bdd_4_lut (.I0(n13745), .I1(n9845), .I2(n13268), .I3(\instruction[11] ), 
            .O(n13748));
    defparam n13745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_12772 (.I0(\instruction[10] ), .I1(n13526), 
            .I2(n11648), .I3(\instruction[11] ), .O(n13745));
    defparam instruction_10__bdd_4_lut_12772.LUT_INIT = 16'he4aa;
    SB_LUT4 n13751_bdd_4_lut (.I0(n13751), .I1(ram_s_13_5), .I2(ram_s_12_5), 
            .I3(\instruction[9] ), .O(n10733));
    defparam n13751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12322 (.I0(\instruction[8] ), .I1(ram_s_14_5), 
            .I2(ram_s_15_5), .I3(\instruction[9] ), .O(n13751));
    defparam instruction_8__bdd_4_lut_12322.LUT_INIT = 16'he4aa;
    SB_LUT4 n13835_bdd_4_lut (.I0(n13835), .I1(ram_s_1_6), .I2(ram_s_0_6), 
            .I3(\instruction[9] ), .O(n13838));
    defparam n13835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12472 (.I0(\instruction[8] ), .I1(ram_s_2_6), 
            .I2(ram_s_3_6), .I3(\instruction[9] ), .O(n13835));
    defparam instruction_8__bdd_4_lut_12472.LUT_INIT = 16'he4aa;
    SB_LUT4 n14015_bdd_4_lut (.I0(n14015), .I1(ram_s_21_7), .I2(ram_s_20_7), 
            .I3(\instruction[9] ), .O(n10355));
    defparam n14015_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12517 (.I0(\instruction[8] ), .I1(ram_s_22_7), 
            .I2(ram_s_23_7), .I3(\instruction[9] ), .O(n14015));
    defparam instruction_8__bdd_4_lut_12517.LUT_INIT = 16'he4aa;
    SB_LUT4 n14069_bdd_4_lut (.I0(n14069), .I1(ram_s_13_4), .I2(ram_s_12_4), 
            .I3(\instruction[9] ), .O(n14072));
    defparam n14069_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12572 (.I0(\instruction[8] ), .I1(ram_s_14_4), 
            .I2(ram_s_15_4), .I3(\instruction[9] ), .O(n14069));
    defparam instruction_8__bdd_4_lut_12572.LUT_INIT = 16'he4aa;
    SB_LUT4 n14135_bdd_4_lut (.I0(n14135), .I1(ram_s_17_6), .I2(ram_s_16_6), 
            .I3(\instruction[9] ), .O(n9560));
    defparam n14135_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12827 (.I0(\instruction[8] ), .I1(ram_s_18_6), 
            .I2(ram_s_19_6), .I3(\instruction[9] ), .O(n14135));
    defparam instruction_8__bdd_4_lut_12827.LUT_INIT = 16'he4aa;
    SB_LUT4 n14375_bdd_4_lut (.I0(n14375), .I1(n13220), .I2(n13838), .I3(\instruction[11] ), 
            .O(n14378));
    defparam n14375_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut_13112 (.I0(\instruction[10] ), .I1(n11306), 
            .I2(n9464), .I3(\instruction[11] ), .O(n14375));
    defparam instruction_10__bdd_4_lut_13112.LUT_INIT = 16'he4aa;
    SB_LUT4 n14441_bdd_4_lut (.I0(n14441), .I1(ram_s_17_7), .I2(ram_s_16_7), 
            .I3(\instruction[9] ), .O(n10310));
    defparam n14441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_12942 (.I0(\instruction[8] ), .I1(ram_s_18_7), 
            .I2(ram_s_19_7), .I3(\instruction[9] ), .O(n14441));
    defparam instruction_8__bdd_4_lut_12942.LUT_INIT = 16'he4aa;
    SB_LUT4 n14579_bdd_4_lut (.I0(n14579), .I1(ram_s_5_4), .I2(ram_s_4_4), 
            .I3(\instruction[9] ), .O(n14582));
    defparam n14579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_13002 (.I0(\instruction[8] ), .I1(ram_s_6_4), 
            .I2(ram_s_7_4), .I3(\instruction[9] ), .O(n14579));
    defparam instruction_8__bdd_4_lut_13002.LUT_INIT = 16'he4aa;
    SB_LUT4 n14651_bdd_4_lut (.I0(n14651), .I1(ram_s_9_5), .I2(ram_s_8_5), 
            .I3(\instruction[9] ), .O(n10643));
    defparam n14651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_13102 (.I0(\instruction[8] ), .I1(ram_s_10_5), 
            .I2(ram_s_11_5), .I3(\instruction[9] ), .O(n14651));
    defparam instruction_8__bdd_4_lut_13102.LUT_INIT = 16'he4aa;
    SB_LUT4 n14771_bdd_4_lut (.I0(n14771), .I1(ram_s_29_5), .I2(ram_s_28_5), 
            .I3(\instruction[9] ), .O(n8948));
    defparam n14771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_13212 (.I0(\instruction[8] ), .I1(ram_s_30_5), 
            .I2(ram_s_31_5), .I3(\instruction[9] ), .O(n14771));
    defparam instruction_8__bdd_4_lut_13212.LUT_INIT = 16'he4aa;
    SB_LUT4 n14783_bdd_4_lut (.I0(n14783), .I1(n14582), .I2(n11522), .I3(\instruction[11] ), 
            .O(n14786));
    defparam n14783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_10__bdd_4_lut (.I0(\instruction[10] ), .I1(n12728), 
            .I2(n14072), .I3(\instruction[11] ), .O(n14783));
    defparam instruction_10__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14903_bdd_4_lut (.I0(n14903), .I1(ram_s_13_7), .I2(ram_s_12_7), 
            .I3(\instruction[9] ), .O(n10262));
    defparam n14903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_13267 (.I0(\instruction[8] ), .I1(ram_s_14_7), 
            .I2(ram_s_15_7), .I3(\instruction[9] ), .O(n14903));
    defparam instruction_8__bdd_4_lut_13267.LUT_INIT = 16'he4aa;
    SB_LUT4 n14969_bdd_4_lut (.I0(n14969), .I1(ram_s_13_6), .I2(ram_s_12_6), 
            .I3(\instruction[9] ), .O(n9464));
    defparam n14969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_13312 (.I0(\instruction[8] ), .I1(ram_s_14_6), 
            .I2(ram_s_15_6), .I3(\instruction[9] ), .O(n14969));
    defparam instruction_8__bdd_4_lut_13312.LUT_INIT = 16'he4aa;
    SB_LUT4 n15023_bdd_4_lut (.I0(n15023), .I1(ram_s_21_4), .I2(ram_s_20_4), 
            .I3(\instruction[9] ), .O(n9845));
    defparam n15023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut_13492 (.I0(\instruction[8] ), .I1(ram_s_22_4), 
            .I2(ram_s_23_4), .I3(\instruction[9] ), .O(n15023));
    defparam instruction_8__bdd_4_lut_13492.LUT_INIT = 16'he4aa;
    SB_LUT4 n15239_bdd_4_lut (.I0(n15239), .I1(ram_s_9_7), .I2(ram_s_8_7), 
            .I3(\instruction[9] ), .O(n10235));
    defparam n15239_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 instruction_8__bdd_4_lut (.I0(\instruction[8] ), .I1(ram_s_10_7), 
            .I2(ram_s_11_7), .I3(\instruction[9] ), .O(n15239));
    defparam instruction_8__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i7767_3_lut (.I0(ram_s_4_2), .I1(ram_s_5_2), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n8826));
    defparam i7767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7768_3_lut (.I0(ram_s_6_2), .I1(ram_s_7_2), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n8827));
    defparam i7768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7750_3_lut (.I0(ram_s_2_2), .I1(ram_s_3_2), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n8809));
    defparam i7750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7749_3_lut (.I0(ram_s_0_2), .I1(ram_s_1_2), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n8808));
    defparam i7749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8598_3_lut (.I0(ram_s_4_3), .I1(ram_s_5_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n9657));
    defparam i8598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8599_3_lut (.I0(ram_s_6_3), .I1(ram_s_7_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n9658));
    defparam i8599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8221_3_lut (.I0(ram_s_2_3), .I1(ram_s_3_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n9280));
    defparam i8221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8220_3_lut (.I0(ram_s_0_3), .I1(ram_s_1_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n9279));
    defparam i8220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7747_3_lut (.I0(n12434), .I1(n13568), .I2(\instruction[10] ), 
            .I3(wea[0]), .O(n8806));
    defparam i7747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7741_3_lut (.I0(n11864), .I1(n11834), .I2(\instruction[10] ), 
            .I3(wea[0]), .O(n8800));
    defparam i7741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10014_3_lut (.I0(ram_s_20_1), .I1(ram_s_21_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11073));
    defparam i10014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10015_3_lut (.I0(ram_s_22_1), .I1(ram_s_23_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11074));
    defparam i10015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10006_3_lut (.I0(ram_s_18_1), .I1(ram_s_19_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11065));
    defparam i10006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10005_3_lut (.I0(ram_s_16_1), .I1(ram_s_17_1), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n11064));
    defparam i10005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i30_2_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n30));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i30_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i33_2_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n33));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i33_2_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i32_2_lut_4_lut (.I0(n7), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n32));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i32_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i35_2_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n35));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i35_2_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i34_2_lut_4_lut (.I0(n6), .I1(\instruction[9] ), 
            .I2(\instruction[10] ), .I3(\instruction[11] ), .O(n34));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i34_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7935_3_lut (.I0(n13724), .I1(n11438), .I2(\instruction[10] ), 
            .I3(wea[0]), .O(n8994));
    defparam i7935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7936_3_lut (.I0(n13742), .I1(n12134), .I2(\instruction[10] ), 
            .I3(wea[0]), .O(n8995));
    defparam i7936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8974_3_lut (.I0(ram_s_10_3), .I1(ram_s_11_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n10033));
    defparam i8974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8973_3_lut (.I0(ram_s_8_3), .I1(ram_s_9_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n10032));
    defparam i8973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9231_3_lut (.I0(ram_s_12_3), .I1(ram_s_13_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n10290));
    defparam i9231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9232_3_lut (.I0(ram_s_14_3), .I1(ram_s_15_3), .I2(\instruction[8] ), 
            .I3(wea[0]), .O(n10291));
    defparam i9232_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module state_machine
//

module state_machine (n8580, bram_enable, CLK_3P3_MHZ_c, \t_state[1] , 
            t_state_2__N_28, internal_reset, BTN1_c, run, \stack_pointer_carry[4] , 
            wea, special_bit, internal_reset_N_50, \instruction[13] , 
            instruction_13_N_701, t_state_1_N_95, loadstar_type, \sy_addr[4] , 
            sx_addr4_value);
    input n8580;
    output bram_enable;
    input CLK_3P3_MHZ_c;
    output \t_state[1] ;
    input t_state_2__N_28;
    output internal_reset;
    input BTN1_c;
    output run;
    input \stack_pointer_carry[4] ;
    input [0:0]wea;
    input special_bit;
    output internal_reset_N_50;
    input \instruction[13] ;
    output instruction_13_N_701;
    output t_state_1_N_95;
    input loadstar_type;
    input \sy_addr[4] ;
    output sx_addr4_value;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    wire n4344, n546, run_value_N_30, n8623;
    
    SB_DFF t_state_i2 (.Q(bram_enable), .C(CLK_3P3_MHZ_c), .D(n8580));   // src/state_machine.vhd(70[9] 79[16])
    SB_DFFSR t_state_i1 (.Q(\t_state[1] ), .C(CLK_3P3_MHZ_c), .D(n4344), 
            .R(t_state_2__N_28));   // src/state_machine.vhd(70[9] 79[16])
    SB_DFFSS internal_reset_117 (.Q(internal_reset), .C(CLK_3P3_MHZ_c), 
            .D(n546), .S(BTN1_c));   // src/state_machine.vhd(70[9] 79[16])
    SB_DFFSS run_116 (.Q(run), .C(CLK_3P3_MHZ_c), .D(run_value_N_30), 
            .S(n8623));   // src/state_machine.vhd(70[9] 79[16])
    SB_LUT4 i1_3_lut (.I0(run), .I1(bram_enable), .I2(\stack_pointer_carry[4] ), 
            .I3(wea[0]), .O(n546));   // src/state_machine.vhd(108[26:84])
    defparam i1_3_lut.LUT_INIT = 16'hd5d5;
    SB_LUT4 i10110_3_lut (.I0(internal_reset), .I1(\t_state[1] ), .I2(special_bit), 
            .I3(wea[0]), .O(n4344));
    defparam i10110_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 internal_reset_I_0_1_lut (.I0(internal_reset), .I1(wea[0]), 
            .I2(wea[0]), .I3(wea[0]), .O(internal_reset_N_50));   // src/state_machine.vhd(123[24:42])
    defparam internal_reset_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(bram_enable), .I1(BTN1_c), .I2(\stack_pointer_carry[4] ), 
            .I3(internal_reset), .O(n8623));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1300;
    SB_LUT4 i1_2_lut_4_lut_adj_299 (.I0(bram_enable), .I1(BTN1_c), .I2(\stack_pointer_carry[4] ), 
            .I3(run), .O(run_value_N_30));
    defparam i1_2_lut_4_lut_adj_299.LUT_INIT = 16'h1300;
    SB_LUT4 instruction_13_I_0_39_1_lut (.I0(\instruction[13] ), .I1(wea[0]), 
            .I2(wea[0]), .I3(wea[0]), .O(instruction_13_N_701));   // src/sel_of_out_port_value.vhd(140[15:33])
    defparam instruction_13_I_0_39_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 t_state_1_I_0_47_1_lut (.I0(\t_state[1] ), .I1(wea[0]), .I2(wea[0]), 
            .I3(wea[0]), .O(t_state_1_N_95));   // src/register_bank_control.vhd(93[17:30])
    defparam t_state_1_I_0_47_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i609_3_lut (.I0(loadstar_type), .I1(\sy_addr[4] ), .I2(bram_enable), 
            .I3(wea[0]), .O(sx_addr4_value));   // src/state_machine.vhd(158[21] 160[56])
    defparam i609_3_lut.LUT_INIT = 16'hc6c6;
    
endmodule
//
// Verilog Description of module stack
//

module stack (CLK_3P3_MHZ_c, shadow_zero_flag, shadow_bank, special_bit, 
            shadow_carry_flag, \stack_pointer_carry[4] , wea, bram_enable, 
            t_state_2__N_28, pop_stack, \t_state[1] , internal_reset, 
            t_state_1_N_95, push_stack_N_165, pop_stack_N_164, \instruction[12] , 
            carry_flag, zero_flag, \sy_addr[4] , run, address, VCC_net, 
            stack_memory);
    input CLK_3P3_MHZ_c;
    output shadow_zero_flag;
    output shadow_bank;
    output special_bit;
    output shadow_carry_flag;
    output \stack_pointer_carry[4] ;
    input [0:0]wea;
    input bram_enable;
    output t_state_2__N_28;
    input pop_stack;
    input \t_state[1] ;
    input internal_reset;
    input t_state_1_N_95;
    input push_stack_N_165;
    input pop_stack_N_164;
    input \instruction[12] ;
    input carry_flag;
    input zero_flag;
    input \sy_addr[4] ;
    input run;
    input [11:0]address;
    input VCC_net;
    output [11:0]stack_memory;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [7:0]data_out_ram_low;   // src/stack.vhd(112[12:28])
    
    wire shadow_zero_value;
    wire [4:0]n12;
    wire [4:0]stack_pointer;   // src/stack.vhd(111[12:25])
    wire [4:0]stack_pointer_carry;   // src/stack.vhd(57[9:28])
    wire [4:0]half_pointer_value;   // src/stack.vhd(120[12:30])
    
    wire n6_adj_884, n4268, stack_pointer_value_0__N_636, n8229, n8651, 
        stack_pointer_value_0__N_609, n249;
    
    SB_DFF shadow_zero_value_160 (.Q(shadow_zero_value), .C(CLK_3P3_MHZ_c), 
           .D(data_out_ram_low[1]));   // src/stack.vhd(130[9] 136[16])
    SB_DFF shadow_zero_flag_161 (.Q(shadow_zero_flag), .C(CLK_3P3_MHZ_c), 
           .D(shadow_zero_value));   // src/stack.vhd(130[9] 136[16])
    SB_DFF shadow_bank_162 (.Q(shadow_bank), .C(CLK_3P3_MHZ_c), .D(data_out_ram_low[2]));   // src/stack.vhd(130[9] 136[16])
    SB_DFF special_bit_163 (.Q(special_bit), .C(CLK_3P3_MHZ_c), .D(data_out_ram_low[3]));   // src/stack.vhd(130[9] 136[16])
    SB_DFF shadow_carry_flag_159 (.Q(shadow_carry_flag), .C(CLK_3P3_MHZ_c), 
           .D(data_out_ram_low[0]));   // src/stack.vhd(130[9] 136[16])
    SB_DFF stack_pointer__i0 (.Q(stack_pointer[0]), .C(CLK_3P3_MHZ_c), .D(n12[0]));   // src/stack.vhd(140[9] 146[16])
    SB_DFF stack_pointer__i1 (.Q(stack_pointer[1]), .C(CLK_3P3_MHZ_c), .D(n12[1]));   // src/stack.vhd(140[9] 146[16])
    SB_DFF stack_pointer__i2 (.Q(stack_pointer[2]), .C(CLK_3P3_MHZ_c), .D(n12[2]));   // src/stack.vhd(140[9] 146[16])
    SB_LUT4 stack_pointer_carry_3__I_0_3_lut (.I0(stack_pointer[4]), .I1(stack_pointer_carry[3]), 
            .I2(half_pointer_value[4]), .I3(wea[0]), .O(\stack_pointer_carry[4] ));   // src/stack.vhd(400[9] 407[18])
    defparam stack_pointer_carry_3__I_0_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 t_state_2__I_0_137_1_lut (.I0(bram_enable), .I1(wea[0]), .I2(wea[0]), 
            .I3(wea[0]), .O(t_state_2__N_28));   // src/state_machine.vhd(123[66:80])
    defparam t_state_2__I_0_137_1_lut.LUT_INIT = 16'h5555;
    SB_DFF stack_pointer__i3 (.Q(stack_pointer[3]), .C(CLK_3P3_MHZ_c), .D(n12[3]));   // src/stack.vhd(140[9] 146[16])
    SB_DFF stack_pointer__i4 (.Q(stack_pointer[4]), .C(CLK_3P3_MHZ_c), .D(n12[4]));   // src/stack.vhd(140[9] 146[16])
    SB_LUT4 i3_4_lut (.I0(stack_pointer[0]), .I1(n6_adj_884), .I2(pop_stack), 
            .I3(n4268), .O(stack_pointer_carry[0]));   // src/stack.vhd(348[9] 355[18])
    defparam i3_4_lut.LUT_INIT = 16'h8808;
    SB_LUT4 i1_2_lut (.I0(\t_state[1] ), .I1(n4268), .I2(wea[0]), .I3(wea[0]), 
            .O(stack_pointer_value_0__N_636));   // src/stack.vhd(247[4:52])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 stack_pointer_carry_0__I_0_3_lut (.I0(stack_pointer[1]), .I1(stack_pointer_carry[0]), 
            .I2(half_pointer_value[1]), .I3(wea[0]), .O(stack_pointer_carry[1]));   // src/stack.vhd(361[9] 368[18])
    defparam stack_pointer_carry_0__I_0_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 stack_pointer_carry_1__I_0_3_lut (.I0(stack_pointer[2]), .I1(stack_pointer_carry[1]), 
            .I2(half_pointer_value[2]), .I3(wea[0]), .O(stack_pointer_carry[2]));   // src/stack.vhd(374[9] 381[18])
    defparam stack_pointer_carry_1__I_0_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 stack_pointer_carry_2__I_0_3_lut (.I0(stack_pointer[3]), .I1(stack_pointer_carry[2]), 
            .I2(half_pointer_value[3]), .I3(wea[0]), .O(stack_pointer_carry[3]));   // src/stack.vhd(387[9] 394[18])
    defparam stack_pointer_carry_2__I_0_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4059_3_lut (.I0(half_pointer_value[4]), .I1(internal_reset), 
            .I2(stack_pointer_carry[3]), .I3(wea[0]), .O(n12[4]));   // src/stack.vhd(140[9] 146[16])
    defparam i4059_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i4058_3_lut (.I0(half_pointer_value[3]), .I1(internal_reset), 
            .I2(stack_pointer_carry[2]), .I3(wea[0]), .O(n12[3]));   // src/stack.vhd(140[9] 146[16])
    defparam i4058_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i4057_3_lut (.I0(half_pointer_value[2]), .I1(internal_reset), 
            .I2(stack_pointer_carry[1]), .I3(wea[0]), .O(n12[2]));   // src/stack.vhd(140[9] 146[16])
    defparam i4057_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i4056_3_lut (.I0(half_pointer_value[1]), .I1(internal_reset), 
            .I2(stack_pointer_carry[0]), .I3(wea[0]), .O(n12[1]));   // src/stack.vhd(140[9] 146[16])
    defparam i4056_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i2_4_lut (.I0(stack_pointer_value_0__N_636), .I1(pop_stack), 
            .I2(bram_enable), .I3(t_state_1_N_95), .O(n8229));   // src/stack.vhd(247[4:95])
    defparam i2_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i2_4_lut_adj_298 (.I0(bram_enable), .I1(n8229), .I2(push_stack_N_165), 
            .I3(t_state_1_N_95), .O(n8651));   // src/stack.vhd(242[3] 247[96])
    defparam i2_4_lut_adj_298.LUT_INIT = 16'hcecc;
    SB_LUT4 i4045_4_lut (.I0(stack_pointer_value_0__N_609), .I1(internal_reset), 
            .I2(stack_pointer[0]), .I3(n8651), .O(n12[0]));   // src/stack.vhd(140[9] 146[16])
    defparam i4045_4_lut.LUT_INIT = 16'h2322;
    SB_LUT4 i2_4_lut_4_lut (.I0(bram_enable), .I1(\t_state[1] ), .I2(stack_pointer[0]), 
            .I3(pop_stack_N_164), .O(stack_pointer_value_0__N_609));   // src/stack.vhd(242[3] 244[73])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h5010;
    SB_LUT4 i607_3_lut_4_lut (.I0(\t_state[1] ), .I1(n4268), .I2(n249), 
            .I3(stack_pointer[4]), .O(half_pointer_value[4]));   // src/stack.vhd(340[3] 343[78])
    defparam i607_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 i606_3_lut_4_lut (.I0(\t_state[1] ), .I1(n4268), .I2(n249), 
            .I3(stack_pointer[3]), .O(half_pointer_value[3]));   // src/stack.vhd(340[3] 343[78])
    defparam i606_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 i605_3_lut_4_lut (.I0(\t_state[1] ), .I1(n4268), .I2(n249), 
            .I3(stack_pointer[2]), .O(half_pointer_value[2]));   // src/stack.vhd(340[3] 343[78])
    defparam i605_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 i603_3_lut_4_lut (.I0(\t_state[1] ), .I1(n4268), .I2(n249), 
            .I3(stack_pointer[1]), .O(half_pointer_value[1]));   // src/stack.vhd(340[3] 343[78])
    defparam i603_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 i4029_2_lut_3_lut (.I0(bram_enable), .I1(pop_stack_N_164), .I2(\instruction[12] ), 
            .I3(wea[0]), .O(n4268));
    defparam i4029_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(bram_enable), .I1(pop_stack_N_164), 
            .I2(\instruction[12] ), .I3(\t_state[1] ), .O(n6_adj_884));
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'hfbaa;
    SB_LUT4 half_pointer_value_4__I_249_i1_2_lut_4_lut_4_lut (.I0(bram_enable), 
            .I1(pop_stack_N_164), .I2(\instruction[12] ), .I3(\t_state[1] ), 
            .O(n249));
    defparam half_pointer_value_4__I_249_i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h04ff;
    \ram(16,5)  stack_ram (.stack_pointer({stack_pointer}), .n12({n12}), 
            .carry_flag(carry_flag), .zero_flag(zero_flag), .\sy_addr[4] (\sy_addr[4] ), 
            .run(run), .address({address}), .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), 
            .\t_state[1] (\t_state[1] ), .VCC_net(VCC_net), .wea({wea}), 
            .stack_memory({stack_memory}), .\data_out_ram_low[3] (data_out_ram_low[3]), 
            .\data_out_ram_low[2] (data_out_ram_low[2]), .\data_out_ram_low[1] (data_out_ram_low[1]), 
            .\data_out_ram_low[0] (data_out_ram_low[0]));   // src/stack.vhd(185[14:17])
    
endmodule
//
// Verilog Description of module \ram(16,5) 
//

module \ram(16,5)  (stack_pointer, n12, carry_flag, zero_flag, \sy_addr[4] , 
            run, address, CLK_3P3_MHZ_c, \t_state[1] , VCC_net, wea, 
            stack_memory, \data_out_ram_low[3] , \data_out_ram_low[2] , 
            \data_out_ram_low[1] , \data_out_ram_low[0] );
    input [4:0]stack_pointer;
    input [4:0]n12;
    input carry_flag;
    input zero_flag;
    input \sy_addr[4] ;
    input run;
    input [11:0]address;
    input CLK_3P3_MHZ_c;
    input \t_state[1] ;
    input VCC_net;
    input [0:0]wea;
    output [11:0]stack_memory;
    output \data_out_ram_low[3] ;
    output \data_out_ram_low[2] ;
    output \data_out_ram_low[1] ;
    output \data_out_ram_low[0] ;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    SB_RAM256x16 ram_s0 (.RDATA({stack_memory, \data_out_ram_low[3] , \data_out_ram_low[2] , 
            \data_out_ram_low[1] , \data_out_ram_low[0] }), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(VCC_net), .RE(VCC_net), .RADDR({wea, wea, wea, 
            n12}), .WCLK(CLK_3P3_MHZ_c), .WCLKE(VCC_net), .WE(\t_state[1] ), 
            .WADDR({wea, wea, wea, stack_pointer}), .MASK({wea, wea, 
            wea, wea, wea, wea, wea, wea, wea, wea, wea, wea, 
            wea, wea, wea, wea}), .WDATA({address, run, \sy_addr[4] , 
            zero_flag, carry_flag}));
    defparam ram_s0.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam ram_s0.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    
endmodule
//
// Verilog Description of module spm_with_output_reg
//

module spm_with_output_reg (spm_data, CLK_3P3_MHZ_c, port_id, ram_s_70_3, 
            ram_s_71_3, ram_s_69_3, ram_s_68_3, \sx[7] , \sx[6] , 
            \sx[5] , \sx[4] , \register_vector[10] , ram_s_34_7, ram_s_35_7, 
            ram_s_33_7, ram_s_32_7, \register_vector[9] , ram_s_11_6, 
            ram_s_8_6, \register_vector[11] , ram_s_62_4, ram_s_63_4, 
            ram_s_2_7, ram_s_3_7, ram_s_1_7, ram_s_0_7, ram_s_66_4, 
            ram_s_67_4, ram_s_65_4, ram_s_64_4, \register_vector[8] , 
            ram_s_142_3, ram_s_141_3, ram_s_140_3, ram_s_209_3, ram_s_130_0, 
            ram_s_131_0, ram_s_129_0, ram_s_128_0, ram_s_70_4, ram_s_71_4, 
            ram_s_69_4, ram_s_68_4, ram_s_171_5, ram_s_168_5, ram_s_14_6, 
            ram_s_13_6, ram_s_12_6, ram_s_202_1, ram_s_203_1, ram_s_6_5, 
            ram_s_7_5, ram_s_14_5, ram_s_5_5, ram_s_4_5, ram_s_13_5, 
            ram_s_12_5, ram_s_43_2, ram_s_2_0, ram_s_3_0, ram_s_2_1, 
            ram_s_3_1, ram_s_1_0, ram_s_0_0, ram_s_66_0, ram_s_67_0, 
            ram_s_34_1, ram_s_35_1, ram_s_33_1, ram_s_32_1, ram_s_201_1, 
            ram_s_200_1, ram_s_1_1, ram_s_0_1, ram_s_65_0, ram_s_64_0, 
            ram_s_11_2, ram_s_8_2, ram_s_38_0, ram_s_39_0, ram_s_40_2, 
            ram_s_74_7, ram_s_75_7, ram_s_73_7, ram_s_72_7, ram_s_130_7, 
            ram_s_131_7, ram_s_129_7, ram_s_128_7, ram_s_37_0, ram_s_36_0, 
            ram_s_142_5, ram_s_141_5, ram_s_140_5, ram_s_62_0, ram_s_63_0, 
            ram_s_194_1, ram_s_195_1, ram_s_193_1, ram_s_192_1, ram_s_74_4, 
            ram_s_75_4, ram_s_73_4, ram_s_72_4, ram_s_43_7, ram_s_40_7, 
            ram_s_74_2, ram_s_75_2, ram_s_73_2, ram_s_72_2, ram_s_186_3, 
            ram_s_185_3, ram_s_190_2, ram_s_191_2, ram_s_43_1, wea, 
            ram_s_40_1, ram_s_6_7, ram_s_7_7, ram_s_134_0, ram_s_135_0, 
            ram_s_5_7, ram_s_4_7, ram_s_133_0, ram_s_132_0, ram_s_34_2, 
            ram_s_35_2, ram_s_58_5, ram_s_58_0, ram_s_57_0, ram_s_139_0, 
            ram_s_136_0, ram_s_190_5, ram_s_191_5, ram_s_57_5, ram_s_33_2, 
            ram_s_32_2, ram_s_142_7, ram_s_141_7, ram_s_140_7, ram_s_81_5, 
            ram_s_190_1, ram_s_191_1, ram_s_139_1, ram_s_136_1, ram_s_38_7, 
            ram_s_39_7, ram_s_37_7, ram_s_36_7, n893, ram_s_14_4, 
            ram_s_190_7, ram_s_191_7, ram_s_47_2, ram_s_45_2, ram_s_44_2, 
            ram_s_134_5, ram_s_135_5, ram_s_133_5, ram_s_132_5, n2567, 
            ram_s_209_7, n2566, ram_s_209_6, n2565, ram_s_209_5, n2564, 
            ram_s_209_4, n2563, n2562, ram_s_209_2, n2561, ram_s_209_1, 
            n2560, ram_s_209_0, n2519, ram_s_203_7, n2518, ram_s_203_6, 
            n2517, ram_s_203_5, n2516, ram_s_203_4, n2515, ram_s_203_3, 
            n2514, ram_s_203_2, n2513, n2512, ram_s_203_0, n2511, 
            ram_s_202_7, n2510, ram_s_202_6, n2509, ram_s_202_5, n2508, 
            ram_s_202_4, n2507, ram_s_202_3, n2506, ram_s_202_2, n2505, 
            n2504, ram_s_202_0, n2503, ram_s_201_7, n2502, ram_s_201_6, 
            n2501, ram_s_201_5, n2500, ram_s_201_4, n2499, ram_s_201_3, 
            n2498, ram_s_201_2, n2497, n2496, ram_s_201_0, n2495, 
            ram_s_200_7, n2494, ram_s_200_6, n2493, ram_s_200_5, n2492, 
            ram_s_200_4, n2491, ram_s_200_3, n2490, ram_s_200_2, n2489, 
            n2488, ram_s_200_0, n2487, ram_s_199_7, n2486, ram_s_199_6, 
            n2485, ram_s_199_5, n2484, ram_s_199_4, n2483, ram_s_199_3, 
            n2482, ram_s_199_2, n2481, ram_s_199_1, n2480, ram_s_199_0, 
            n2479, ram_s_198_7, n2478, ram_s_198_6, n2477, ram_s_198_5, 
            n2476, ram_s_198_4, n2475, ram_s_198_3, n2474, ram_s_198_2, 
            n2473, ram_s_198_1, n2472, ram_s_198_0, n2471, ram_s_197_7, 
            n2470, ram_s_197_6, n2469, ram_s_197_5, n2468, ram_s_197_4, 
            n2467, ram_s_197_3, n2466, ram_s_197_2, n2465, ram_s_197_1, 
            n2464, ram_s_197_0, n2463, ram_s_196_7, n2462, ram_s_196_6, 
            n2461, ram_s_196_5, n2460, ram_s_196_4, n2459, ram_s_196_3, 
            n2458, ram_s_196_2, n2457, ram_s_196_1, n2456, ram_s_196_0, 
            n2455, ram_s_195_7, n2454, ram_s_195_6, n2453, ram_s_195_5, 
            n2452, ram_s_195_4, n2451, ram_s_195_3, n2450, ram_s_195_2, 
            n2449, n2448, ram_s_195_0, n2447, ram_s_194_7, n2446, 
            ram_s_194_6, n2445, ram_s_194_5, n2444, ram_s_194_4, n2443, 
            ram_s_194_3, n2442, ram_s_194_2, n2441, n2440, ram_s_194_0, 
            n2439, ram_s_193_7, n2438, ram_s_193_6, n2437, ram_s_193_5, 
            n2436, ram_s_193_4, n2435, ram_s_193_3, n2434, ram_s_193_2, 
            n2433, n2432, ram_s_193_0, n2431, ram_s_192_7, n2430, 
            ram_s_192_6, n2429, ram_s_192_5, n2428, ram_s_192_4, n2427, 
            ram_s_192_3, n2426, ram_s_192_2, n2425, n2424, ram_s_192_0, 
            n2423, n2422, ram_s_191_6, n2421, n2420, ram_s_191_4, 
            n2419, ram_s_191_3, n2418, n2417, n2416, ram_s_191_0, 
            n2415, n2414, ram_s_190_6, n2413, n2412, ram_s_190_4, 
            n2411, ram_s_190_3, n2410, n2409, n2408, ram_s_190_0, 
            n2383, ram_s_186_7, n2382, ram_s_186_6, n2381, ram_s_186_5, 
            n2380, ram_s_186_4, n2379, n2378, ram_s_186_2, n2377, 
            ram_s_186_1, n2376, ram_s_186_0, n2375, ram_s_185_7, n2374, 
            ram_s_185_6, n2373, ram_s_185_5, n2372, ram_s_185_4, n2371, 
            n2370, ram_s_185_2, n2369, ram_s_185_1, n2368, ram_s_185_0, 
            n2295, ram_s_175_7, n2294, ram_s_175_6, n2293, ram_s_175_5, 
            n2292, ram_s_175_4, n2291, ram_s_175_3, n2290, ram_s_175_2, 
            n2289, ram_s_175_1, n2288, ram_s_175_0, n2279, ram_s_173_7, 
            n2278, ram_s_173_6, n2277, ram_s_173_5, n2276, ram_s_173_4, 
            n2275, ram_s_173_3, n2274, ram_s_173_2, n2273, ram_s_173_1, 
            n2272, ram_s_173_0, n2271, ram_s_172_7, n2270, ram_s_172_6, 
            n2269, ram_s_172_5, n2268, ram_s_172_4, n2267, ram_s_172_3, 
            n2266, ram_s_172_2, n2265, ram_s_172_1, n2264, ram_s_172_0, 
            n2263, ram_s_171_7, n2262, ram_s_171_6, n2261, n2260, 
            ram_s_171_4, n2259, ram_s_171_3, n2258, ram_s_171_2, n2257, 
            ram_s_171_1, n2256, ram_s_171_0, n2239, ram_s_168_7, n2238, 
            ram_s_168_6, n2237, n2236, ram_s_168_4, n2235, ram_s_168_3, 
            n2234, ram_s_168_2, n2233, ram_s_168_1, n2232, ram_s_168_0, 
            n2231, ram_s_167_7, n2230, ram_s_167_6, n2229, ram_s_167_5, 
            n2228, ram_s_167_4, n2227, ram_s_167_3, n2226, ram_s_167_2, 
            n2225, ram_s_167_1, n2224, ram_s_167_0, n2223, ram_s_166_7, 
            n2222, ram_s_166_6, n2221, ram_s_166_5, n2220, ram_s_166_4, 
            n2219, ram_s_166_3, n2218, ram_s_166_2, n2217, ram_s_166_1, 
            n2216, ram_s_166_0, n2215, ram_s_165_7, n2214, ram_s_165_6, 
            n2213, ram_s_165_5, n2212, ram_s_165_4, n2211, ram_s_165_3, 
            n2210, ram_s_165_2, n2209, ram_s_165_1, n2208, ram_s_165_0, 
            n2207, ram_s_164_7, n2206, ram_s_164_6, n2205, ram_s_164_5, 
            n2204, ram_s_164_4, n2203, ram_s_164_3, n2202, ram_s_164_2, 
            n2201, ram_s_164_1, n2200, ram_s_164_0, n2199, ram_s_163_7, 
            n2198, ram_s_163_6, n2197, ram_s_163_5, n2196, ram_s_163_4, 
            n2195, ram_s_163_3, n2194, ram_s_163_2, n2193, ram_s_163_1, 
            n2192, ram_s_163_0, n2191, ram_s_162_7, n2190, ram_s_162_6, 
            n2189, ram_s_162_5, n2188, ram_s_162_4, n2187, ram_s_162_3, 
            n2186, ram_s_162_2, n2185, ram_s_162_1, n2184, ram_s_162_0, 
            n2183, ram_s_161_7, n2182, ram_s_161_6, n2181, ram_s_161_5, 
            n2180, ram_s_161_4, n2179, ram_s_161_3, n2178, ram_s_161_2, 
            n2177, ram_s_161_1, n2176, ram_s_161_0, n2175, ram_s_160_7, 
            n2174, ram_s_160_6, n2173, ram_s_160_5, n2172, ram_s_160_4, 
            n2171, ram_s_160_3, n2170, ram_s_160_2, n2169, ram_s_160_1, 
            n2168, ram_s_160_0, n2031, n2030, ram_s_142_6, n2029, 
            n2028, ram_s_142_4, n2027, n2026, ram_s_142_2, n2025, 
            ram_s_142_1, n2024, ram_s_142_0, n2023, n2022, ram_s_141_6, 
            n2021, n2020, ram_s_141_4, n2019, n2018, ram_s_141_2, 
            n2017, ram_s_141_1, n2016, ram_s_141_0, n2015, n2014, 
            ram_s_140_6, n2013, n2012, ram_s_140_4, n2011, n2010, 
            ram_s_140_2, n2009, ram_s_140_1, n2008, ram_s_140_0, n2007, 
            ram_s_139_7, n2006, ram_s_139_6, n2005, ram_s_139_5, n2004, 
            ram_s_139_4, n2003, ram_s_139_3, n2002, ram_s_139_2, n2001, 
            n2000, n1983, ram_s_136_7, n1982, ram_s_136_6, n1981, 
            ram_s_136_5, n1980, ram_s_136_4, n1979, ram_s_136_3, n1978, 
            ram_s_136_2, n1977, n1976, n1975, ram_s_135_7, n1974, 
            ram_s_135_6, n1973, n1972, ram_s_135_4, n1971, ram_s_135_3, 
            n1970, ram_s_135_2, n1969, ram_s_135_1, n1968, n1967, 
            ram_s_134_7, n1966, ram_s_134_6, n1965, n1964, ram_s_134_4, 
            n1963, ram_s_134_3, n1962, ram_s_134_2, n1961, ram_s_134_1, 
            n1960, n1959, ram_s_133_7, n1958, ram_s_133_6, n1957, 
            n1956, ram_s_133_4, n1955, ram_s_133_3, n1954, ram_s_133_2, 
            n1953, ram_s_133_1, n1952, n1951, ram_s_132_7, n1950, 
            ram_s_132_6, n1949, n1948, ram_s_132_4, n1947, ram_s_132_3, 
            n1946, ram_s_132_2, n1945, ram_s_132_1, n1944, n1943, 
            n1942, ram_s_131_6, n1941, ram_s_131_5, n1940, ram_s_131_4, 
            n1939, ram_s_131_3, n1938, ram_s_131_2, n1937, ram_s_131_1, 
            n1936, n1935, n1934, ram_s_130_6, n1933, ram_s_130_5, 
            n1932, ram_s_130_4, n1931, ram_s_130_3, n1930, ram_s_130_2, 
            n1929, ram_s_130_1, n1928, n1927, n1926, ram_s_129_6, 
            n1925, ram_s_129_5, n1924, ram_s_129_4, n1923, ram_s_129_3, 
            n1922, ram_s_129_2, n1921, ram_s_129_1, n1920, n1919, 
            n1918, ram_s_128_6, n1917, ram_s_128_5, n1916, ram_s_128_4, 
            n1915, ram_s_128_3, n1914, ram_s_128_2, n1913, ram_s_128_1, 
            n1912, n1543, ram_s_81_7, n1542, ram_s_81_6, n1541, 
            n1540, ram_s_81_4, n1539, ram_s_81_3, n1538, ram_s_81_2, 
            n1537, ram_s_81_1, n1536, ram_s_81_0, n1495, n1494, 
            ram_s_75_6, n1493, ram_s_75_5, n1492, n1491, ram_s_75_3, 
            n1490, n1489, ram_s_75_1, n1488, ram_s_75_0, n1487, 
            n1486, ram_s_74_6, n1485, ram_s_74_5, n1484, n1483, 
            ram_s_74_3, n1482, n1481, ram_s_74_1, n1480, ram_s_74_0, 
            n1479, n1478, ram_s_73_6, n1477, ram_s_73_5, n1476, 
            n1475, ram_s_73_3, n1474, n1473, ram_s_73_1, n1472, 
            ram_s_73_0, n1471, n1470, ram_s_72_6, n1469, ram_s_72_5, 
            n1468, n1467, ram_s_72_3, n1466, n1465, ram_s_72_1, 
            n1464, ram_s_72_0, n1463, ram_s_71_7, n1462, ram_s_71_6, 
            n1461, ram_s_71_5, n1460, n1459, n1458, ram_s_71_2, 
            n1457, ram_s_71_1, n1456, ram_s_71_0, n1455, ram_s_70_7, 
            n1454, ram_s_70_6, n1453, ram_s_70_5, n1452, n1451, 
            n1450, ram_s_70_2, n1449, ram_s_70_1, n1448, ram_s_70_0, 
            n1447, ram_s_69_7, n1446, ram_s_69_6, n1445, ram_s_69_5, 
            n1444, n1443, n1442, ram_s_69_2, n1441, ram_s_69_1, 
            n1440, ram_s_69_0, n1439, ram_s_68_7, n1438, ram_s_68_6, 
            n1437, ram_s_68_5, n1436, n1435, n1434, ram_s_68_2, 
            n1433, ram_s_68_1, n1432, ram_s_68_0, n1431, ram_s_67_7, 
            n1430, ram_s_67_6, n1429, ram_s_67_5, n1428, n1427, 
            ram_s_67_3, n1426, ram_s_67_2, n1425, ram_s_67_1, n1424, 
            n1423, ram_s_66_7, n1422, ram_s_66_6, n1421, ram_s_66_5, 
            n1420, n1419, ram_s_66_3, n1418, ram_s_66_2, n1417, 
            ram_s_66_1, n1416, n1415, ram_s_65_7, n1414, ram_s_65_6, 
            n1413, ram_s_65_5, n1412, n1411, ram_s_65_3, n1410, 
            ram_s_65_2, n1409, ram_s_65_1, n1408, n1407, ram_s_64_7, 
            n1406, ram_s_64_6, n1405, ram_s_64_5, n1404, n1403, 
            ram_s_64_3, n1402, ram_s_64_2, n1401, ram_s_64_1, n1400, 
            n1399, ram_s_63_7, n1398, ram_s_63_6, n1397, ram_s_63_5, 
            n1396, n1395, ram_s_63_3, n1394, ram_s_63_2, n1393, 
            ram_s_63_1, n1392, n1391, ram_s_62_7, n1390, ram_s_62_6, 
            n1389, ram_s_62_5, n1388, n1387, ram_s_62_3, n1386, 
            ram_s_62_2, n1385, ram_s_62_1, n1384, n1359, ram_s_58_7, 
            n1358, ram_s_58_6, n1357, n1356, ram_s_58_4, n1355, 
            ram_s_58_3, n1354, ram_s_58_2, n1353, ram_s_58_1, n1352, 
            n1351, ram_s_57_7, n1350, ram_s_57_6, n1349, n1348, 
            ram_s_57_4, n1347, ram_s_57_3, n1346, ram_s_57_2, n1345, 
            ram_s_57_1, n1344, n1271, ram_s_47_7, n1270, ram_s_47_6, 
            n1269, ram_s_47_5, n1268, ram_s_47_4, n1267, ram_s_47_3, 
            n1266, n1265, ram_s_47_1, n1264, ram_s_47_0, n1255, 
            ram_s_45_7, n1254, ram_s_45_6, n1253, ram_s_45_5, n1252, 
            ram_s_45_4, n1251, ram_s_45_3, n1250, n1249, ram_s_45_1, 
            n1248, ram_s_45_0, n1247, ram_s_44_7, n1246, ram_s_44_6, 
            n1245, ram_s_44_5, n1244, ram_s_44_4, n1243, ram_s_44_3, 
            n1242, n1241, ram_s_44_1, n1240, ram_s_44_0, n1239, 
            n1238, ram_s_43_6, n1237, ram_s_43_5, n1236, ram_s_43_4, 
            n1235, ram_s_43_3, n1234, n1233, n1232, ram_s_43_0, 
            n1215, n1214, ram_s_40_6, n1213, ram_s_40_5, n1212, 
            ram_s_40_4, n1211, ram_s_40_3, n1210, n1209, n1208, 
            ram_s_40_0, n1207, n1206, ram_s_39_6, n1205, ram_s_39_5, 
            n1204, ram_s_39_4, n1203, ram_s_39_3, n1202, ram_s_39_2, 
            n1201, ram_s_39_1, n1200, n1199, n1198, ram_s_38_6, 
            n1197, ram_s_38_5, n1196, ram_s_38_4, n1195, ram_s_38_3, 
            n1194, ram_s_38_2, n1193, ram_s_38_1, n1192, n1191, 
            n1190, ram_s_37_6, n1189, ram_s_37_5, n1188, ram_s_37_4, 
            n1187, ram_s_37_3, n1186, ram_s_37_2, n1185, ram_s_37_1, 
            n1184, n1183, n1182, ram_s_36_6, n1181, ram_s_36_5, 
            n1180, ram_s_36_4, n1179, ram_s_36_3, n1178, ram_s_36_2, 
            n1177, ram_s_36_1, n1176, n1175, n1174, ram_s_35_6, 
            n1173, ram_s_35_5, n1172, ram_s_35_4, n1171, ram_s_35_3, 
            n1170, n1169, n1168, ram_s_35_0, n1167, n1166, ram_s_34_6, 
            n1165, ram_s_34_5, n1164, ram_s_34_4, n1163, ram_s_34_3, 
            n1162, n1161, n1160, ram_s_34_0, n1159, n1158, ram_s_33_6, 
            n1157, ram_s_33_5, n1156, ram_s_33_4, n1155, ram_s_33_3, 
            n1154, n1153, n1152, ram_s_33_0, n1151, n1150, ram_s_32_6, 
            n1149, ram_s_32_5, n1148, ram_s_32_4, n1147, ram_s_32_3, 
            n1146, n1145, n1144, ram_s_32_0, n1051, n1047, n1046, 
            n1045, ram_s_0_2, n1044, ram_s_12_3, n1043, n1042, ram_s_11_1, 
            n1041, n1040, ram_s_12_1, n1038, ram_s_11_4, n182, n1037, 
            ram_s_12_4, n54, n1036, ram_s_11_7, n183, n1035, n55, 
            n1034, ram_s_12_7, n184, n1033, ram_s_12_2, n56, n1032, 
            ram_s_11_5, n185, n1031, n57, n1030, ram_s_12_0, n186, 
            n1029, ram_s_11_3, n58, n187, n59, n188, n60, n189, 
            n61, n190, n62, n191, n63, n192, n1017, ram_s_0_3, 
            n64, n1016, ram_s_0_4, n193, n1015, ram_s_0_5, n65, 
            n1014, ram_s_0_6, n194, n1013, n66, n1012, n195, n1011, 
            n67, n1010, ram_s_1_2, n1009, ram_s_1_3, n1008, ram_s_1_4, 
            n1007, ram_s_1_5, n1006, ram_s_4_4, n1005, n1004, n1003, 
            ram_s_5_0, n1002, ram_s_4_6, n1001, ram_s_5_1, n998, 
            ram_s_8_5, n997, n996, n995, ram_s_7_4, n994, ram_s_7_1, 
            n993, ram_s_6_6, n992, ram_s_6_3, n989, n988, ram_s_8_3, 
            n987, ram_s_8_0, n986, n199, n985, ram_s_7_2, n71, 
            n984, n200, n983, ram_s_6_4, n72, n980, ram_s_8_7, 
            n979, ram_s_8_4, n978, ram_s_8_1, n977, ram_s_7_6, n976, 
            ram_s_7_3, n975, ram_s_7_0, n974, n973, ram_s_1_6, n972, 
            n971, n970, n969, ram_s_2_2, n968, ram_s_2_3, n967, 
            ram_s_2_4, n966, ram_s_2_5, n965, ram_s_2_6, n964, n963, 
            n962, n961, ram_s_3_2, n960, ram_s_3_3, n959, ram_s_3_4, 
            n958, ram_s_3_5, n957, ram_s_14_7, n952, ram_s_3_6, 
            n950, n946, ram_s_4_0, n944, ram_s_4_1, n941, ram_s_4_2, 
            n940, ram_s_5_2, n939, ram_s_5_3, n935, n934, ram_s_6_0, 
            n933, ram_s_6_1, n932, ram_s_6_2, n931, ram_s_5_6, n930, 
            n927, ram_s_4_3, n926, n925, ram_s_13_3, n924, ram_s_13_4, 
            n923, n210, n82, n212, n84, n213, n85, n214, n86, 
            n217, n89, n218, n90, n219, n91, n220, n92, n221, 
            n93, n222, n94, n223, n95, n224, n96, n225, n97, 
            n918, ram_s_13_7, n917, ram_s_14_0, n916, ram_s_14_1, 
            spm_enable, n244, n116, n115, n243, n245, n117, n246, 
            n118, n48, n176, n249, n121, n250, n122, n251, n123, 
            n252, n124, n253, n125, n254, n126, n255, n127, 
            n256, n128, n257, n129, ram_s_14_2, ram_s_13_2, ram_s_11_0, 
            n911, n909, n908, ram_s_14_3, n907, ram_s_13_1, n906, 
            n904, ram_s_13_0, n901, ram_s_5_4, n899);
    output [7:0]spm_data;
    input CLK_3P3_MHZ_c;
    input [7:0]port_id;
    output ram_s_70_3;
    output ram_s_71_3;
    output ram_s_69_3;
    output ram_s_68_3;
    input \sx[7] ;
    input \sx[6] ;
    input \sx[5] ;
    input \sx[4] ;
    input \register_vector[10] ;
    output ram_s_34_7;
    output ram_s_35_7;
    output ram_s_33_7;
    output ram_s_32_7;
    input \register_vector[9] ;
    output ram_s_11_6;
    output ram_s_8_6;
    input \register_vector[11] ;
    output ram_s_62_4;
    output ram_s_63_4;
    output ram_s_2_7;
    output ram_s_3_7;
    output ram_s_1_7;
    output ram_s_0_7;
    output ram_s_66_4;
    output ram_s_67_4;
    output ram_s_65_4;
    output ram_s_64_4;
    input \register_vector[8] ;
    output ram_s_142_3;
    output ram_s_141_3;
    output ram_s_140_3;
    output ram_s_209_3;
    output ram_s_130_0;
    output ram_s_131_0;
    output ram_s_129_0;
    output ram_s_128_0;
    output ram_s_70_4;
    output ram_s_71_4;
    output ram_s_69_4;
    output ram_s_68_4;
    output ram_s_171_5;
    output ram_s_168_5;
    output ram_s_14_6;
    output ram_s_13_6;
    output ram_s_12_6;
    output ram_s_202_1;
    output ram_s_203_1;
    output ram_s_6_5;
    output ram_s_7_5;
    output ram_s_14_5;
    output ram_s_5_5;
    output ram_s_4_5;
    output ram_s_13_5;
    output ram_s_12_5;
    output ram_s_43_2;
    output ram_s_2_0;
    output ram_s_3_0;
    output ram_s_2_1;
    output ram_s_3_1;
    output ram_s_1_0;
    output ram_s_0_0;
    output ram_s_66_0;
    output ram_s_67_0;
    output ram_s_34_1;
    output ram_s_35_1;
    output ram_s_33_1;
    output ram_s_32_1;
    output ram_s_201_1;
    output ram_s_200_1;
    output ram_s_1_1;
    output ram_s_0_1;
    output ram_s_65_0;
    output ram_s_64_0;
    output ram_s_11_2;
    output ram_s_8_2;
    output ram_s_38_0;
    output ram_s_39_0;
    output ram_s_40_2;
    output ram_s_74_7;
    output ram_s_75_7;
    output ram_s_73_7;
    output ram_s_72_7;
    output ram_s_130_7;
    output ram_s_131_7;
    output ram_s_129_7;
    output ram_s_128_7;
    output ram_s_37_0;
    output ram_s_36_0;
    output ram_s_142_5;
    output ram_s_141_5;
    output ram_s_140_5;
    output ram_s_62_0;
    output ram_s_63_0;
    output ram_s_194_1;
    output ram_s_195_1;
    output ram_s_193_1;
    output ram_s_192_1;
    output ram_s_74_4;
    output ram_s_75_4;
    output ram_s_73_4;
    output ram_s_72_4;
    output ram_s_43_7;
    output ram_s_40_7;
    output ram_s_74_2;
    output ram_s_75_2;
    output ram_s_73_2;
    output ram_s_72_2;
    output ram_s_186_3;
    output ram_s_185_3;
    output ram_s_190_2;
    output ram_s_191_2;
    output ram_s_43_1;
    input [0:0]wea;
    output ram_s_40_1;
    output ram_s_6_7;
    output ram_s_7_7;
    output ram_s_134_0;
    output ram_s_135_0;
    output ram_s_5_7;
    output ram_s_4_7;
    output ram_s_133_0;
    output ram_s_132_0;
    output ram_s_34_2;
    output ram_s_35_2;
    output ram_s_58_5;
    output ram_s_58_0;
    output ram_s_57_0;
    output ram_s_139_0;
    output ram_s_136_0;
    output ram_s_190_5;
    output ram_s_191_5;
    output ram_s_57_5;
    output ram_s_33_2;
    output ram_s_32_2;
    output ram_s_142_7;
    output ram_s_141_7;
    output ram_s_140_7;
    output ram_s_81_5;
    output ram_s_190_1;
    output ram_s_191_1;
    output ram_s_139_1;
    output ram_s_136_1;
    output ram_s_38_7;
    output ram_s_39_7;
    output ram_s_37_7;
    output ram_s_36_7;
    input n893;
    output ram_s_14_4;
    output ram_s_190_7;
    output ram_s_191_7;
    output ram_s_47_2;
    output ram_s_45_2;
    output ram_s_44_2;
    output ram_s_134_5;
    output ram_s_135_5;
    output ram_s_133_5;
    output ram_s_132_5;
    input n2567;
    output ram_s_209_7;
    input n2566;
    output ram_s_209_6;
    input n2565;
    output ram_s_209_5;
    input n2564;
    output ram_s_209_4;
    input n2563;
    input n2562;
    output ram_s_209_2;
    input n2561;
    output ram_s_209_1;
    input n2560;
    output ram_s_209_0;
    input n2519;
    output ram_s_203_7;
    input n2518;
    output ram_s_203_6;
    input n2517;
    output ram_s_203_5;
    input n2516;
    output ram_s_203_4;
    input n2515;
    output ram_s_203_3;
    input n2514;
    output ram_s_203_2;
    input n2513;
    input n2512;
    output ram_s_203_0;
    input n2511;
    output ram_s_202_7;
    input n2510;
    output ram_s_202_6;
    input n2509;
    output ram_s_202_5;
    input n2508;
    output ram_s_202_4;
    input n2507;
    output ram_s_202_3;
    input n2506;
    output ram_s_202_2;
    input n2505;
    input n2504;
    output ram_s_202_0;
    input n2503;
    output ram_s_201_7;
    input n2502;
    output ram_s_201_6;
    input n2501;
    output ram_s_201_5;
    input n2500;
    output ram_s_201_4;
    input n2499;
    output ram_s_201_3;
    input n2498;
    output ram_s_201_2;
    input n2497;
    input n2496;
    output ram_s_201_0;
    input n2495;
    output ram_s_200_7;
    input n2494;
    output ram_s_200_6;
    input n2493;
    output ram_s_200_5;
    input n2492;
    output ram_s_200_4;
    input n2491;
    output ram_s_200_3;
    input n2490;
    output ram_s_200_2;
    input n2489;
    input n2488;
    output ram_s_200_0;
    input n2487;
    output ram_s_199_7;
    input n2486;
    output ram_s_199_6;
    input n2485;
    output ram_s_199_5;
    input n2484;
    output ram_s_199_4;
    input n2483;
    output ram_s_199_3;
    input n2482;
    output ram_s_199_2;
    input n2481;
    output ram_s_199_1;
    input n2480;
    output ram_s_199_0;
    input n2479;
    output ram_s_198_7;
    input n2478;
    output ram_s_198_6;
    input n2477;
    output ram_s_198_5;
    input n2476;
    output ram_s_198_4;
    input n2475;
    output ram_s_198_3;
    input n2474;
    output ram_s_198_2;
    input n2473;
    output ram_s_198_1;
    input n2472;
    output ram_s_198_0;
    input n2471;
    output ram_s_197_7;
    input n2470;
    output ram_s_197_6;
    input n2469;
    output ram_s_197_5;
    input n2468;
    output ram_s_197_4;
    input n2467;
    output ram_s_197_3;
    input n2466;
    output ram_s_197_2;
    input n2465;
    output ram_s_197_1;
    input n2464;
    output ram_s_197_0;
    input n2463;
    output ram_s_196_7;
    input n2462;
    output ram_s_196_6;
    input n2461;
    output ram_s_196_5;
    input n2460;
    output ram_s_196_4;
    input n2459;
    output ram_s_196_3;
    input n2458;
    output ram_s_196_2;
    input n2457;
    output ram_s_196_1;
    input n2456;
    output ram_s_196_0;
    input n2455;
    output ram_s_195_7;
    input n2454;
    output ram_s_195_6;
    input n2453;
    output ram_s_195_5;
    input n2452;
    output ram_s_195_4;
    input n2451;
    output ram_s_195_3;
    input n2450;
    output ram_s_195_2;
    input n2449;
    input n2448;
    output ram_s_195_0;
    input n2447;
    output ram_s_194_7;
    input n2446;
    output ram_s_194_6;
    input n2445;
    output ram_s_194_5;
    input n2444;
    output ram_s_194_4;
    input n2443;
    output ram_s_194_3;
    input n2442;
    output ram_s_194_2;
    input n2441;
    input n2440;
    output ram_s_194_0;
    input n2439;
    output ram_s_193_7;
    input n2438;
    output ram_s_193_6;
    input n2437;
    output ram_s_193_5;
    input n2436;
    output ram_s_193_4;
    input n2435;
    output ram_s_193_3;
    input n2434;
    output ram_s_193_2;
    input n2433;
    input n2432;
    output ram_s_193_0;
    input n2431;
    output ram_s_192_7;
    input n2430;
    output ram_s_192_6;
    input n2429;
    output ram_s_192_5;
    input n2428;
    output ram_s_192_4;
    input n2427;
    output ram_s_192_3;
    input n2426;
    output ram_s_192_2;
    input n2425;
    input n2424;
    output ram_s_192_0;
    input n2423;
    input n2422;
    output ram_s_191_6;
    input n2421;
    input n2420;
    output ram_s_191_4;
    input n2419;
    output ram_s_191_3;
    input n2418;
    input n2417;
    input n2416;
    output ram_s_191_0;
    input n2415;
    input n2414;
    output ram_s_190_6;
    input n2413;
    input n2412;
    output ram_s_190_4;
    input n2411;
    output ram_s_190_3;
    input n2410;
    input n2409;
    input n2408;
    output ram_s_190_0;
    input n2383;
    output ram_s_186_7;
    input n2382;
    output ram_s_186_6;
    input n2381;
    output ram_s_186_5;
    input n2380;
    output ram_s_186_4;
    input n2379;
    input n2378;
    output ram_s_186_2;
    input n2377;
    output ram_s_186_1;
    input n2376;
    output ram_s_186_0;
    input n2375;
    output ram_s_185_7;
    input n2374;
    output ram_s_185_6;
    input n2373;
    output ram_s_185_5;
    input n2372;
    output ram_s_185_4;
    input n2371;
    input n2370;
    output ram_s_185_2;
    input n2369;
    output ram_s_185_1;
    input n2368;
    output ram_s_185_0;
    input n2295;
    output ram_s_175_7;
    input n2294;
    output ram_s_175_6;
    input n2293;
    output ram_s_175_5;
    input n2292;
    output ram_s_175_4;
    input n2291;
    output ram_s_175_3;
    input n2290;
    output ram_s_175_2;
    input n2289;
    output ram_s_175_1;
    input n2288;
    output ram_s_175_0;
    input n2279;
    output ram_s_173_7;
    input n2278;
    output ram_s_173_6;
    input n2277;
    output ram_s_173_5;
    input n2276;
    output ram_s_173_4;
    input n2275;
    output ram_s_173_3;
    input n2274;
    output ram_s_173_2;
    input n2273;
    output ram_s_173_1;
    input n2272;
    output ram_s_173_0;
    input n2271;
    output ram_s_172_7;
    input n2270;
    output ram_s_172_6;
    input n2269;
    output ram_s_172_5;
    input n2268;
    output ram_s_172_4;
    input n2267;
    output ram_s_172_3;
    input n2266;
    output ram_s_172_2;
    input n2265;
    output ram_s_172_1;
    input n2264;
    output ram_s_172_0;
    input n2263;
    output ram_s_171_7;
    input n2262;
    output ram_s_171_6;
    input n2261;
    input n2260;
    output ram_s_171_4;
    input n2259;
    output ram_s_171_3;
    input n2258;
    output ram_s_171_2;
    input n2257;
    output ram_s_171_1;
    input n2256;
    output ram_s_171_0;
    input n2239;
    output ram_s_168_7;
    input n2238;
    output ram_s_168_6;
    input n2237;
    input n2236;
    output ram_s_168_4;
    input n2235;
    output ram_s_168_3;
    input n2234;
    output ram_s_168_2;
    input n2233;
    output ram_s_168_1;
    input n2232;
    output ram_s_168_0;
    input n2231;
    output ram_s_167_7;
    input n2230;
    output ram_s_167_6;
    input n2229;
    output ram_s_167_5;
    input n2228;
    output ram_s_167_4;
    input n2227;
    output ram_s_167_3;
    input n2226;
    output ram_s_167_2;
    input n2225;
    output ram_s_167_1;
    input n2224;
    output ram_s_167_0;
    input n2223;
    output ram_s_166_7;
    input n2222;
    output ram_s_166_6;
    input n2221;
    output ram_s_166_5;
    input n2220;
    output ram_s_166_4;
    input n2219;
    output ram_s_166_3;
    input n2218;
    output ram_s_166_2;
    input n2217;
    output ram_s_166_1;
    input n2216;
    output ram_s_166_0;
    input n2215;
    output ram_s_165_7;
    input n2214;
    output ram_s_165_6;
    input n2213;
    output ram_s_165_5;
    input n2212;
    output ram_s_165_4;
    input n2211;
    output ram_s_165_3;
    input n2210;
    output ram_s_165_2;
    input n2209;
    output ram_s_165_1;
    input n2208;
    output ram_s_165_0;
    input n2207;
    output ram_s_164_7;
    input n2206;
    output ram_s_164_6;
    input n2205;
    output ram_s_164_5;
    input n2204;
    output ram_s_164_4;
    input n2203;
    output ram_s_164_3;
    input n2202;
    output ram_s_164_2;
    input n2201;
    output ram_s_164_1;
    input n2200;
    output ram_s_164_0;
    input n2199;
    output ram_s_163_7;
    input n2198;
    output ram_s_163_6;
    input n2197;
    output ram_s_163_5;
    input n2196;
    output ram_s_163_4;
    input n2195;
    output ram_s_163_3;
    input n2194;
    output ram_s_163_2;
    input n2193;
    output ram_s_163_1;
    input n2192;
    output ram_s_163_0;
    input n2191;
    output ram_s_162_7;
    input n2190;
    output ram_s_162_6;
    input n2189;
    output ram_s_162_5;
    input n2188;
    output ram_s_162_4;
    input n2187;
    output ram_s_162_3;
    input n2186;
    output ram_s_162_2;
    input n2185;
    output ram_s_162_1;
    input n2184;
    output ram_s_162_0;
    input n2183;
    output ram_s_161_7;
    input n2182;
    output ram_s_161_6;
    input n2181;
    output ram_s_161_5;
    input n2180;
    output ram_s_161_4;
    input n2179;
    output ram_s_161_3;
    input n2178;
    output ram_s_161_2;
    input n2177;
    output ram_s_161_1;
    input n2176;
    output ram_s_161_0;
    input n2175;
    output ram_s_160_7;
    input n2174;
    output ram_s_160_6;
    input n2173;
    output ram_s_160_5;
    input n2172;
    output ram_s_160_4;
    input n2171;
    output ram_s_160_3;
    input n2170;
    output ram_s_160_2;
    input n2169;
    output ram_s_160_1;
    input n2168;
    output ram_s_160_0;
    input n2031;
    input n2030;
    output ram_s_142_6;
    input n2029;
    input n2028;
    output ram_s_142_4;
    input n2027;
    input n2026;
    output ram_s_142_2;
    input n2025;
    output ram_s_142_1;
    input n2024;
    output ram_s_142_0;
    input n2023;
    input n2022;
    output ram_s_141_6;
    input n2021;
    input n2020;
    output ram_s_141_4;
    input n2019;
    input n2018;
    output ram_s_141_2;
    input n2017;
    output ram_s_141_1;
    input n2016;
    output ram_s_141_0;
    input n2015;
    input n2014;
    output ram_s_140_6;
    input n2013;
    input n2012;
    output ram_s_140_4;
    input n2011;
    input n2010;
    output ram_s_140_2;
    input n2009;
    output ram_s_140_1;
    input n2008;
    output ram_s_140_0;
    input n2007;
    output ram_s_139_7;
    input n2006;
    output ram_s_139_6;
    input n2005;
    output ram_s_139_5;
    input n2004;
    output ram_s_139_4;
    input n2003;
    output ram_s_139_3;
    input n2002;
    output ram_s_139_2;
    input n2001;
    input n2000;
    input n1983;
    output ram_s_136_7;
    input n1982;
    output ram_s_136_6;
    input n1981;
    output ram_s_136_5;
    input n1980;
    output ram_s_136_4;
    input n1979;
    output ram_s_136_3;
    input n1978;
    output ram_s_136_2;
    input n1977;
    input n1976;
    input n1975;
    output ram_s_135_7;
    input n1974;
    output ram_s_135_6;
    input n1973;
    input n1972;
    output ram_s_135_4;
    input n1971;
    output ram_s_135_3;
    input n1970;
    output ram_s_135_2;
    input n1969;
    output ram_s_135_1;
    input n1968;
    input n1967;
    output ram_s_134_7;
    input n1966;
    output ram_s_134_6;
    input n1965;
    input n1964;
    output ram_s_134_4;
    input n1963;
    output ram_s_134_3;
    input n1962;
    output ram_s_134_2;
    input n1961;
    output ram_s_134_1;
    input n1960;
    input n1959;
    output ram_s_133_7;
    input n1958;
    output ram_s_133_6;
    input n1957;
    input n1956;
    output ram_s_133_4;
    input n1955;
    output ram_s_133_3;
    input n1954;
    output ram_s_133_2;
    input n1953;
    output ram_s_133_1;
    input n1952;
    input n1951;
    output ram_s_132_7;
    input n1950;
    output ram_s_132_6;
    input n1949;
    input n1948;
    output ram_s_132_4;
    input n1947;
    output ram_s_132_3;
    input n1946;
    output ram_s_132_2;
    input n1945;
    output ram_s_132_1;
    input n1944;
    input n1943;
    input n1942;
    output ram_s_131_6;
    input n1941;
    output ram_s_131_5;
    input n1940;
    output ram_s_131_4;
    input n1939;
    output ram_s_131_3;
    input n1938;
    output ram_s_131_2;
    input n1937;
    output ram_s_131_1;
    input n1936;
    input n1935;
    input n1934;
    output ram_s_130_6;
    input n1933;
    output ram_s_130_5;
    input n1932;
    output ram_s_130_4;
    input n1931;
    output ram_s_130_3;
    input n1930;
    output ram_s_130_2;
    input n1929;
    output ram_s_130_1;
    input n1928;
    input n1927;
    input n1926;
    output ram_s_129_6;
    input n1925;
    output ram_s_129_5;
    input n1924;
    output ram_s_129_4;
    input n1923;
    output ram_s_129_3;
    input n1922;
    output ram_s_129_2;
    input n1921;
    output ram_s_129_1;
    input n1920;
    input n1919;
    input n1918;
    output ram_s_128_6;
    input n1917;
    output ram_s_128_5;
    input n1916;
    output ram_s_128_4;
    input n1915;
    output ram_s_128_3;
    input n1914;
    output ram_s_128_2;
    input n1913;
    output ram_s_128_1;
    input n1912;
    input n1543;
    output ram_s_81_7;
    input n1542;
    output ram_s_81_6;
    input n1541;
    input n1540;
    output ram_s_81_4;
    input n1539;
    output ram_s_81_3;
    input n1538;
    output ram_s_81_2;
    input n1537;
    output ram_s_81_1;
    input n1536;
    output ram_s_81_0;
    input n1495;
    input n1494;
    output ram_s_75_6;
    input n1493;
    output ram_s_75_5;
    input n1492;
    input n1491;
    output ram_s_75_3;
    input n1490;
    input n1489;
    output ram_s_75_1;
    input n1488;
    output ram_s_75_0;
    input n1487;
    input n1486;
    output ram_s_74_6;
    input n1485;
    output ram_s_74_5;
    input n1484;
    input n1483;
    output ram_s_74_3;
    input n1482;
    input n1481;
    output ram_s_74_1;
    input n1480;
    output ram_s_74_0;
    input n1479;
    input n1478;
    output ram_s_73_6;
    input n1477;
    output ram_s_73_5;
    input n1476;
    input n1475;
    output ram_s_73_3;
    input n1474;
    input n1473;
    output ram_s_73_1;
    input n1472;
    output ram_s_73_0;
    input n1471;
    input n1470;
    output ram_s_72_6;
    input n1469;
    output ram_s_72_5;
    input n1468;
    input n1467;
    output ram_s_72_3;
    input n1466;
    input n1465;
    output ram_s_72_1;
    input n1464;
    output ram_s_72_0;
    input n1463;
    output ram_s_71_7;
    input n1462;
    output ram_s_71_6;
    input n1461;
    output ram_s_71_5;
    input n1460;
    input n1459;
    input n1458;
    output ram_s_71_2;
    input n1457;
    output ram_s_71_1;
    input n1456;
    output ram_s_71_0;
    input n1455;
    output ram_s_70_7;
    input n1454;
    output ram_s_70_6;
    input n1453;
    output ram_s_70_5;
    input n1452;
    input n1451;
    input n1450;
    output ram_s_70_2;
    input n1449;
    output ram_s_70_1;
    input n1448;
    output ram_s_70_0;
    input n1447;
    output ram_s_69_7;
    input n1446;
    output ram_s_69_6;
    input n1445;
    output ram_s_69_5;
    input n1444;
    input n1443;
    input n1442;
    output ram_s_69_2;
    input n1441;
    output ram_s_69_1;
    input n1440;
    output ram_s_69_0;
    input n1439;
    output ram_s_68_7;
    input n1438;
    output ram_s_68_6;
    input n1437;
    output ram_s_68_5;
    input n1436;
    input n1435;
    input n1434;
    output ram_s_68_2;
    input n1433;
    output ram_s_68_1;
    input n1432;
    output ram_s_68_0;
    input n1431;
    output ram_s_67_7;
    input n1430;
    output ram_s_67_6;
    input n1429;
    output ram_s_67_5;
    input n1428;
    input n1427;
    output ram_s_67_3;
    input n1426;
    output ram_s_67_2;
    input n1425;
    output ram_s_67_1;
    input n1424;
    input n1423;
    output ram_s_66_7;
    input n1422;
    output ram_s_66_6;
    input n1421;
    output ram_s_66_5;
    input n1420;
    input n1419;
    output ram_s_66_3;
    input n1418;
    output ram_s_66_2;
    input n1417;
    output ram_s_66_1;
    input n1416;
    input n1415;
    output ram_s_65_7;
    input n1414;
    output ram_s_65_6;
    input n1413;
    output ram_s_65_5;
    input n1412;
    input n1411;
    output ram_s_65_3;
    input n1410;
    output ram_s_65_2;
    input n1409;
    output ram_s_65_1;
    input n1408;
    input n1407;
    output ram_s_64_7;
    input n1406;
    output ram_s_64_6;
    input n1405;
    output ram_s_64_5;
    input n1404;
    input n1403;
    output ram_s_64_3;
    input n1402;
    output ram_s_64_2;
    input n1401;
    output ram_s_64_1;
    input n1400;
    input n1399;
    output ram_s_63_7;
    input n1398;
    output ram_s_63_6;
    input n1397;
    output ram_s_63_5;
    input n1396;
    input n1395;
    output ram_s_63_3;
    input n1394;
    output ram_s_63_2;
    input n1393;
    output ram_s_63_1;
    input n1392;
    input n1391;
    output ram_s_62_7;
    input n1390;
    output ram_s_62_6;
    input n1389;
    output ram_s_62_5;
    input n1388;
    input n1387;
    output ram_s_62_3;
    input n1386;
    output ram_s_62_2;
    input n1385;
    output ram_s_62_1;
    input n1384;
    input n1359;
    output ram_s_58_7;
    input n1358;
    output ram_s_58_6;
    input n1357;
    input n1356;
    output ram_s_58_4;
    input n1355;
    output ram_s_58_3;
    input n1354;
    output ram_s_58_2;
    input n1353;
    output ram_s_58_1;
    input n1352;
    input n1351;
    output ram_s_57_7;
    input n1350;
    output ram_s_57_6;
    input n1349;
    input n1348;
    output ram_s_57_4;
    input n1347;
    output ram_s_57_3;
    input n1346;
    output ram_s_57_2;
    input n1345;
    output ram_s_57_1;
    input n1344;
    input n1271;
    output ram_s_47_7;
    input n1270;
    output ram_s_47_6;
    input n1269;
    output ram_s_47_5;
    input n1268;
    output ram_s_47_4;
    input n1267;
    output ram_s_47_3;
    input n1266;
    input n1265;
    output ram_s_47_1;
    input n1264;
    output ram_s_47_0;
    input n1255;
    output ram_s_45_7;
    input n1254;
    output ram_s_45_6;
    input n1253;
    output ram_s_45_5;
    input n1252;
    output ram_s_45_4;
    input n1251;
    output ram_s_45_3;
    input n1250;
    input n1249;
    output ram_s_45_1;
    input n1248;
    output ram_s_45_0;
    input n1247;
    output ram_s_44_7;
    input n1246;
    output ram_s_44_6;
    input n1245;
    output ram_s_44_5;
    input n1244;
    output ram_s_44_4;
    input n1243;
    output ram_s_44_3;
    input n1242;
    input n1241;
    output ram_s_44_1;
    input n1240;
    output ram_s_44_0;
    input n1239;
    input n1238;
    output ram_s_43_6;
    input n1237;
    output ram_s_43_5;
    input n1236;
    output ram_s_43_4;
    input n1235;
    output ram_s_43_3;
    input n1234;
    input n1233;
    input n1232;
    output ram_s_43_0;
    input n1215;
    input n1214;
    output ram_s_40_6;
    input n1213;
    output ram_s_40_5;
    input n1212;
    output ram_s_40_4;
    input n1211;
    output ram_s_40_3;
    input n1210;
    input n1209;
    input n1208;
    output ram_s_40_0;
    input n1207;
    input n1206;
    output ram_s_39_6;
    input n1205;
    output ram_s_39_5;
    input n1204;
    output ram_s_39_4;
    input n1203;
    output ram_s_39_3;
    input n1202;
    output ram_s_39_2;
    input n1201;
    output ram_s_39_1;
    input n1200;
    input n1199;
    input n1198;
    output ram_s_38_6;
    input n1197;
    output ram_s_38_5;
    input n1196;
    output ram_s_38_4;
    input n1195;
    output ram_s_38_3;
    input n1194;
    output ram_s_38_2;
    input n1193;
    output ram_s_38_1;
    input n1192;
    input n1191;
    input n1190;
    output ram_s_37_6;
    input n1189;
    output ram_s_37_5;
    input n1188;
    output ram_s_37_4;
    input n1187;
    output ram_s_37_3;
    input n1186;
    output ram_s_37_2;
    input n1185;
    output ram_s_37_1;
    input n1184;
    input n1183;
    input n1182;
    output ram_s_36_6;
    input n1181;
    output ram_s_36_5;
    input n1180;
    output ram_s_36_4;
    input n1179;
    output ram_s_36_3;
    input n1178;
    output ram_s_36_2;
    input n1177;
    output ram_s_36_1;
    input n1176;
    input n1175;
    input n1174;
    output ram_s_35_6;
    input n1173;
    output ram_s_35_5;
    input n1172;
    output ram_s_35_4;
    input n1171;
    output ram_s_35_3;
    input n1170;
    input n1169;
    input n1168;
    output ram_s_35_0;
    input n1167;
    input n1166;
    output ram_s_34_6;
    input n1165;
    output ram_s_34_5;
    input n1164;
    output ram_s_34_4;
    input n1163;
    output ram_s_34_3;
    input n1162;
    input n1161;
    input n1160;
    output ram_s_34_0;
    input n1159;
    input n1158;
    output ram_s_33_6;
    input n1157;
    output ram_s_33_5;
    input n1156;
    output ram_s_33_4;
    input n1155;
    output ram_s_33_3;
    input n1154;
    input n1153;
    input n1152;
    output ram_s_33_0;
    input n1151;
    input n1150;
    output ram_s_32_6;
    input n1149;
    output ram_s_32_5;
    input n1148;
    output ram_s_32_4;
    input n1147;
    output ram_s_32_3;
    input n1146;
    input n1145;
    input n1144;
    output ram_s_32_0;
    input n1051;
    input n1047;
    input n1046;
    input n1045;
    output ram_s_0_2;
    input n1044;
    output ram_s_12_3;
    input n1043;
    input n1042;
    output ram_s_11_1;
    input n1041;
    input n1040;
    output ram_s_12_1;
    input n1038;
    output ram_s_11_4;
    output n182;
    input n1037;
    output ram_s_12_4;
    output n54;
    input n1036;
    output ram_s_11_7;
    output n183;
    input n1035;
    output n55;
    input n1034;
    output ram_s_12_7;
    output n184;
    input n1033;
    output ram_s_12_2;
    output n56;
    input n1032;
    output ram_s_11_5;
    output n185;
    input n1031;
    output n57;
    input n1030;
    output ram_s_12_0;
    output n186;
    input n1029;
    output ram_s_11_3;
    output n58;
    output n187;
    output n59;
    output n188;
    output n60;
    output n189;
    output n61;
    output n190;
    output n62;
    output n191;
    output n63;
    output n192;
    input n1017;
    output ram_s_0_3;
    output n64;
    input n1016;
    output ram_s_0_4;
    output n193;
    input n1015;
    output ram_s_0_5;
    output n65;
    input n1014;
    output ram_s_0_6;
    output n194;
    input n1013;
    output n66;
    input n1012;
    output n195;
    input n1011;
    output n67;
    input n1010;
    output ram_s_1_2;
    input n1009;
    output ram_s_1_3;
    input n1008;
    output ram_s_1_4;
    input n1007;
    output ram_s_1_5;
    input n1006;
    output ram_s_4_4;
    input n1005;
    input n1004;
    input n1003;
    output ram_s_5_0;
    input n1002;
    output ram_s_4_6;
    input n1001;
    output ram_s_5_1;
    input n998;
    output ram_s_8_5;
    input n997;
    input n996;
    input n995;
    output ram_s_7_4;
    input n994;
    output ram_s_7_1;
    input n993;
    output ram_s_6_6;
    input n992;
    output ram_s_6_3;
    input n989;
    input n988;
    output ram_s_8_3;
    input n987;
    output ram_s_8_0;
    input n986;
    output n199;
    input n985;
    output ram_s_7_2;
    output n71;
    input n984;
    output n200;
    input n983;
    output ram_s_6_4;
    output n72;
    input n980;
    output ram_s_8_7;
    input n979;
    output ram_s_8_4;
    input n978;
    output ram_s_8_1;
    input n977;
    output ram_s_7_6;
    input n976;
    output ram_s_7_3;
    input n975;
    output ram_s_7_0;
    input n974;
    input n973;
    output ram_s_1_6;
    input n972;
    input n971;
    input n970;
    input n969;
    output ram_s_2_2;
    input n968;
    output ram_s_2_3;
    input n967;
    output ram_s_2_4;
    input n966;
    output ram_s_2_5;
    input n965;
    output ram_s_2_6;
    input n964;
    input n963;
    input n962;
    input n961;
    output ram_s_3_2;
    input n960;
    output ram_s_3_3;
    input n959;
    output ram_s_3_4;
    input n958;
    output ram_s_3_5;
    input n957;
    output ram_s_14_7;
    input n952;
    output ram_s_3_6;
    input n950;
    input n946;
    output ram_s_4_0;
    input n944;
    output ram_s_4_1;
    input n941;
    output ram_s_4_2;
    input n940;
    output ram_s_5_2;
    input n939;
    output ram_s_5_3;
    input n935;
    input n934;
    output ram_s_6_0;
    input n933;
    output ram_s_6_1;
    input n932;
    output ram_s_6_2;
    input n931;
    output ram_s_5_6;
    input n930;
    input n927;
    output ram_s_4_3;
    input n926;
    input n925;
    output ram_s_13_3;
    input n924;
    output ram_s_13_4;
    input n923;
    output n210;
    output n82;
    output n212;
    output n84;
    output n213;
    output n85;
    output n214;
    output n86;
    output n217;
    output n89;
    output n218;
    output n90;
    output n219;
    output n91;
    output n220;
    output n92;
    output n221;
    output n93;
    output n222;
    output n94;
    output n223;
    output n95;
    output n224;
    output n96;
    output n225;
    output n97;
    input n918;
    output ram_s_13_7;
    input n917;
    output ram_s_14_0;
    input n916;
    output ram_s_14_1;
    input spm_enable;
    output n244;
    output n116;
    output n115;
    output n243;
    output n245;
    output n117;
    output n246;
    output n118;
    output n48;
    output n176;
    output n249;
    output n121;
    output n250;
    output n122;
    output n251;
    output n123;
    output n252;
    output n124;
    output n253;
    output n125;
    output n254;
    output n126;
    output n255;
    output n127;
    output n256;
    output n128;
    output n257;
    output n129;
    output ram_s_14_2;
    output ram_s_13_2;
    output ram_s_11_0;
    input n911;
    input n909;
    input n908;
    output ram_s_14_3;
    input n907;
    output ram_s_13_1;
    input n906;
    input n904;
    output ram_s_13_0;
    input n901;
    output ram_s_5_4;
    input n899;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [7:0]spm_ram_data;   // src/spm_with_output_reg.vhd(99[12:24])
    
    SB_DFF spm_data_i0 (.Q(spm_data[0]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[0]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    SB_DFF spm_data_i1 (.Q(spm_data[1]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[1]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    SB_DFF spm_data_i2 (.Q(spm_data[2]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[2]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    SB_DFF spm_data_i3 (.Q(spm_data[3]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[3]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    SB_DFF spm_data_i4 (.Q(spm_data[4]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[4]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    SB_DFF spm_data_i5 (.Q(spm_data[5]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[5]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    SB_DFF spm_data_i6 (.Q(spm_data[6]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[6]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    SB_DFF spm_data_i7 (.Q(spm_data[7]), .C(CLK_3P3_MHZ_c), .D(spm_ram_data[7]));   // src/spm_with_output_reg.vhd(106[5] 108[12])
    \ram(8,8)  spm_ram (.port_id({port_id}), .ram_s_70_3(ram_s_70_3), .ram_s_71_3(ram_s_71_3), 
            .ram_s_69_3(ram_s_69_3), .ram_s_68_3(ram_s_68_3), .\sx[7] (\sx[7] ), 
            .\sx[6] (\sx[6] ), .\sx[5] (\sx[5] ), .\sx[4] (\sx[4] ), .\register_vector[10] (\register_vector[10] ), 
            .ram_s_34_7(ram_s_34_7), .ram_s_35_7(ram_s_35_7), .ram_s_33_7(ram_s_33_7), 
            .ram_s_32_7(ram_s_32_7), .\register_vector[9] (\register_vector[9] ), 
            .ram_s_11_6(ram_s_11_6), .ram_s_8_6(ram_s_8_6), .\register_vector[11] (\register_vector[11] ), 
            .ram_s_62_4(ram_s_62_4), .ram_s_63_4(ram_s_63_4), .ram_s_2_7(ram_s_2_7), 
            .ram_s_3_7(ram_s_3_7), .ram_s_1_7(ram_s_1_7), .ram_s_0_7(ram_s_0_7), 
            .ram_s_66_4(ram_s_66_4), .ram_s_67_4(ram_s_67_4), .ram_s_65_4(ram_s_65_4), 
            .ram_s_64_4(ram_s_64_4), .\register_vector[8] (\register_vector[8] ), 
            .ram_s_142_3(ram_s_142_3), .ram_s_141_3(ram_s_141_3), .ram_s_140_3(ram_s_140_3), 
            .CLK_3P3_MHZ_c(CLK_3P3_MHZ_c), .ram_s_209_3(ram_s_209_3), .ram_s_130_0(ram_s_130_0), 
            .ram_s_131_0(ram_s_131_0), .ram_s_129_0(ram_s_129_0), .ram_s_128_0(ram_s_128_0), 
            .ram_s_70_4(ram_s_70_4), .ram_s_71_4(ram_s_71_4), .ram_s_69_4(ram_s_69_4), 
            .ram_s_68_4(ram_s_68_4), .ram_s_171_5(ram_s_171_5), .ram_s_168_5(ram_s_168_5), 
            .ram_s_14_6(ram_s_14_6), .ram_s_13_6(ram_s_13_6), .ram_s_12_6(ram_s_12_6), 
            .ram_s_202_1(ram_s_202_1), .ram_s_203_1(ram_s_203_1), .ram_s_6_5(ram_s_6_5), 
            .ram_s_7_5(ram_s_7_5), .ram_s_14_5(ram_s_14_5), .ram_s_5_5(ram_s_5_5), 
            .ram_s_4_5(ram_s_4_5), .ram_s_13_5(ram_s_13_5), .ram_s_12_5(ram_s_12_5), 
            .ram_s_43_2(ram_s_43_2), .ram_s_2_0(ram_s_2_0), .ram_s_3_0(ram_s_3_0), 
            .ram_s_2_1(ram_s_2_1), .ram_s_3_1(ram_s_3_1), .ram_s_1_0(ram_s_1_0), 
            .ram_s_0_0(ram_s_0_0), .ram_s_66_0(ram_s_66_0), .ram_s_67_0(ram_s_67_0), 
            .ram_s_34_1(ram_s_34_1), .ram_s_35_1(ram_s_35_1), .ram_s_33_1(ram_s_33_1), 
            .ram_s_32_1(ram_s_32_1), .ram_s_201_1(ram_s_201_1), .ram_s_200_1(ram_s_200_1), 
            .ram_s_1_1(ram_s_1_1), .ram_s_0_1(ram_s_0_1), .ram_s_65_0(ram_s_65_0), 
            .ram_s_64_0(ram_s_64_0), .ram_s_11_2(ram_s_11_2), .ram_s_8_2(ram_s_8_2), 
            .ram_s_38_0(ram_s_38_0), .ram_s_39_0(ram_s_39_0), .ram_s_40_2(ram_s_40_2), 
            .ram_s_74_7(ram_s_74_7), .ram_s_75_7(ram_s_75_7), .ram_s_73_7(ram_s_73_7), 
            .ram_s_72_7(ram_s_72_7), .ram_s_130_7(ram_s_130_7), .ram_s_131_7(ram_s_131_7), 
            .ram_s_129_7(ram_s_129_7), .ram_s_128_7(ram_s_128_7), .ram_s_37_0(ram_s_37_0), 
            .ram_s_36_0(ram_s_36_0), .ram_s_142_5(ram_s_142_5), .ram_s_141_5(ram_s_141_5), 
            .ram_s_140_5(ram_s_140_5), .ram_s_62_0(ram_s_62_0), .ram_s_63_0(ram_s_63_0), 
            .ram_s_194_1(ram_s_194_1), .ram_s_195_1(ram_s_195_1), .ram_s_193_1(ram_s_193_1), 
            .ram_s_192_1(ram_s_192_1), .ram_s_74_4(ram_s_74_4), .ram_s_75_4(ram_s_75_4), 
            .ram_s_73_4(ram_s_73_4), .ram_s_72_4(ram_s_72_4), .ram_s_43_7(ram_s_43_7), 
            .ram_s_40_7(ram_s_40_7), .ram_s_74_2(ram_s_74_2), .ram_s_75_2(ram_s_75_2), 
            .ram_s_73_2(ram_s_73_2), .ram_s_72_2(ram_s_72_2), .ram_s_186_3(ram_s_186_3), 
            .ram_s_185_3(ram_s_185_3), .ram_s_190_2(ram_s_190_2), .ram_s_191_2(ram_s_191_2), 
            .ram_s_43_1(ram_s_43_1), .wea({wea}), .ram_s_40_1(ram_s_40_1), 
            .ram_s_6_7(ram_s_6_7), .ram_s_7_7(ram_s_7_7), .ram_s_134_0(ram_s_134_0), 
            .ram_s_135_0(ram_s_135_0), .ram_s_5_7(ram_s_5_7), .ram_s_4_7(ram_s_4_7), 
            .ram_s_133_0(ram_s_133_0), .ram_s_132_0(ram_s_132_0), .ram_s_34_2(ram_s_34_2), 
            .ram_s_35_2(ram_s_35_2), .ram_s_58_5(ram_s_58_5), .ram_s_58_0(ram_s_58_0), 
            .ram_s_57_0(ram_s_57_0), .ram_s_139_0(ram_s_139_0), .ram_s_136_0(ram_s_136_0), 
            .ram_s_190_5(ram_s_190_5), .ram_s_191_5(ram_s_191_5), .ram_s_57_5(ram_s_57_5), 
            .ram_s_33_2(ram_s_33_2), .ram_s_32_2(ram_s_32_2), .ram_s_142_7(ram_s_142_7), 
            .ram_s_141_7(ram_s_141_7), .ram_s_140_7(ram_s_140_7), .ram_s_81_5(ram_s_81_5), 
            .ram_s_190_1(ram_s_190_1), .ram_s_191_1(ram_s_191_1), .ram_s_139_1(ram_s_139_1), 
            .ram_s_136_1(ram_s_136_1), .ram_s_38_7(ram_s_38_7), .ram_s_39_7(ram_s_39_7), 
            .ram_s_37_7(ram_s_37_7), .ram_s_36_7(ram_s_36_7), .n893(n893), 
            .ram_s_14_4(ram_s_14_4), .ram_s_190_7(ram_s_190_7), .ram_s_191_7(ram_s_191_7), 
            .ram_s_47_2(ram_s_47_2), .spm_ram_data({spm_ram_data}), .ram_s_45_2(ram_s_45_2), 
            .ram_s_44_2(ram_s_44_2), .ram_s_134_5(ram_s_134_5), .ram_s_135_5(ram_s_135_5), 
            .ram_s_133_5(ram_s_133_5), .ram_s_132_5(ram_s_132_5), .n2567(n2567), 
            .ram_s_209_7(ram_s_209_7), .n2566(n2566), .ram_s_209_6(ram_s_209_6), 
            .n2565(n2565), .ram_s_209_5(ram_s_209_5), .n2564(n2564), .ram_s_209_4(ram_s_209_4), 
            .n2563(n2563), .n2562(n2562), .ram_s_209_2(ram_s_209_2), .n2561(n2561), 
            .ram_s_209_1(ram_s_209_1), .n2560(n2560), .ram_s_209_0(ram_s_209_0), 
            .n2519(n2519), .ram_s_203_7(ram_s_203_7), .n2518(n2518), .ram_s_203_6(ram_s_203_6), 
            .n2517(n2517), .ram_s_203_5(ram_s_203_5), .n2516(n2516), .ram_s_203_4(ram_s_203_4), 
            .n2515(n2515), .ram_s_203_3(ram_s_203_3), .n2514(n2514), .ram_s_203_2(ram_s_203_2), 
            .n2513(n2513), .n2512(n2512), .ram_s_203_0(ram_s_203_0), .n2511(n2511), 
            .ram_s_202_7(ram_s_202_7), .n2510(n2510), .ram_s_202_6(ram_s_202_6), 
            .n2509(n2509), .ram_s_202_5(ram_s_202_5), .n2508(n2508), .ram_s_202_4(ram_s_202_4), 
            .n2507(n2507), .ram_s_202_3(ram_s_202_3), .n2506(n2506), .ram_s_202_2(ram_s_202_2), 
            .n2505(n2505), .n2504(n2504), .ram_s_202_0(ram_s_202_0), .n2503(n2503), 
            .ram_s_201_7(ram_s_201_7), .n2502(n2502), .ram_s_201_6(ram_s_201_6), 
            .n2501(n2501), .ram_s_201_5(ram_s_201_5), .n2500(n2500), .ram_s_201_4(ram_s_201_4), 
            .n2499(n2499), .ram_s_201_3(ram_s_201_3), .n2498(n2498), .ram_s_201_2(ram_s_201_2), 
            .n2497(n2497), .n2496(n2496), .ram_s_201_0(ram_s_201_0), .n2495(n2495), 
            .ram_s_200_7(ram_s_200_7), .n2494(n2494), .ram_s_200_6(ram_s_200_6), 
            .n2493(n2493), .ram_s_200_5(ram_s_200_5), .n2492(n2492), .ram_s_200_4(ram_s_200_4), 
            .n2491(n2491), .ram_s_200_3(ram_s_200_3), .n2490(n2490), .ram_s_200_2(ram_s_200_2), 
            .n2489(n2489), .n2488(n2488), .ram_s_200_0(ram_s_200_0), .n2487(n2487), 
            .ram_s_199_7(ram_s_199_7), .n2486(n2486), .ram_s_199_6(ram_s_199_6), 
            .n2485(n2485), .ram_s_199_5(ram_s_199_5), .n2484(n2484), .ram_s_199_4(ram_s_199_4), 
            .n2483(n2483), .ram_s_199_3(ram_s_199_3), .n2482(n2482), .ram_s_199_2(ram_s_199_2), 
            .n2481(n2481), .ram_s_199_1(ram_s_199_1), .n2480(n2480), .ram_s_199_0(ram_s_199_0), 
            .n2479(n2479), .ram_s_198_7(ram_s_198_7), .n2478(n2478), .ram_s_198_6(ram_s_198_6), 
            .n2477(n2477), .ram_s_198_5(ram_s_198_5), .n2476(n2476), .ram_s_198_4(ram_s_198_4), 
            .n2475(n2475), .ram_s_198_3(ram_s_198_3), .n2474(n2474), .ram_s_198_2(ram_s_198_2), 
            .n2473(n2473), .ram_s_198_1(ram_s_198_1), .n2472(n2472), .ram_s_198_0(ram_s_198_0), 
            .n2471(n2471), .ram_s_197_7(ram_s_197_7), .n2470(n2470), .ram_s_197_6(ram_s_197_6), 
            .n2469(n2469), .ram_s_197_5(ram_s_197_5), .n2468(n2468), .ram_s_197_4(ram_s_197_4), 
            .n2467(n2467), .ram_s_197_3(ram_s_197_3), .n2466(n2466), .ram_s_197_2(ram_s_197_2), 
            .n2465(n2465), .ram_s_197_1(ram_s_197_1), .n2464(n2464), .ram_s_197_0(ram_s_197_0), 
            .n2463(n2463), .ram_s_196_7(ram_s_196_7), .n2462(n2462), .ram_s_196_6(ram_s_196_6), 
            .n2461(n2461), .ram_s_196_5(ram_s_196_5), .n2460(n2460), .ram_s_196_4(ram_s_196_4), 
            .n2459(n2459), .ram_s_196_3(ram_s_196_3), .n2458(n2458), .ram_s_196_2(ram_s_196_2), 
            .n2457(n2457), .ram_s_196_1(ram_s_196_1), .n2456(n2456), .ram_s_196_0(ram_s_196_0), 
            .n2455(n2455), .ram_s_195_7(ram_s_195_7), .n2454(n2454), .ram_s_195_6(ram_s_195_6), 
            .n2453(n2453), .ram_s_195_5(ram_s_195_5), .n2452(n2452), .ram_s_195_4(ram_s_195_4), 
            .n2451(n2451), .ram_s_195_3(ram_s_195_3), .n2450(n2450), .ram_s_195_2(ram_s_195_2), 
            .n2449(n2449), .n2448(n2448), .ram_s_195_0(ram_s_195_0), .n2447(n2447), 
            .ram_s_194_7(ram_s_194_7), .n2446(n2446), .ram_s_194_6(ram_s_194_6), 
            .n2445(n2445), .ram_s_194_5(ram_s_194_5), .n2444(n2444), .ram_s_194_4(ram_s_194_4), 
            .n2443(n2443), .ram_s_194_3(ram_s_194_3), .n2442(n2442), .ram_s_194_2(ram_s_194_2), 
            .n2441(n2441), .n2440(n2440), .ram_s_194_0(ram_s_194_0), .n2439(n2439), 
            .ram_s_193_7(ram_s_193_7), .n2438(n2438), .ram_s_193_6(ram_s_193_6), 
            .n2437(n2437), .ram_s_193_5(ram_s_193_5), .n2436(n2436), .ram_s_193_4(ram_s_193_4), 
            .n2435(n2435), .ram_s_193_3(ram_s_193_3), .n2434(n2434), .ram_s_193_2(ram_s_193_2), 
            .n2433(n2433), .n2432(n2432), .ram_s_193_0(ram_s_193_0), .n2431(n2431), 
            .ram_s_192_7(ram_s_192_7), .n2430(n2430), .ram_s_192_6(ram_s_192_6), 
            .n2429(n2429), .ram_s_192_5(ram_s_192_5), .n2428(n2428), .ram_s_192_4(ram_s_192_4), 
            .n2427(n2427), .ram_s_192_3(ram_s_192_3), .n2426(n2426), .ram_s_192_2(ram_s_192_2), 
            .n2425(n2425), .n2424(n2424), .ram_s_192_0(ram_s_192_0), .n2423(n2423), 
            .n2422(n2422), .ram_s_191_6(ram_s_191_6), .n2421(n2421), .n2420(n2420), 
            .ram_s_191_4(ram_s_191_4), .n2419(n2419), .ram_s_191_3(ram_s_191_3), 
            .n2418(n2418), .n2417(n2417), .n2416(n2416), .ram_s_191_0(ram_s_191_0), 
            .n2415(n2415), .n2414(n2414), .ram_s_190_6(ram_s_190_6), .n2413(n2413), 
            .n2412(n2412), .ram_s_190_4(ram_s_190_4), .n2411(n2411), .ram_s_190_3(ram_s_190_3), 
            .n2410(n2410), .n2409(n2409), .n2408(n2408), .ram_s_190_0(ram_s_190_0), 
            .n2383(n2383), .ram_s_186_7(ram_s_186_7), .n2382(n2382), .ram_s_186_6(ram_s_186_6), 
            .n2381(n2381), .ram_s_186_5(ram_s_186_5), .n2380(n2380), .ram_s_186_4(ram_s_186_4), 
            .n2379(n2379), .n2378(n2378), .ram_s_186_2(ram_s_186_2), .n2377(n2377), 
            .ram_s_186_1(ram_s_186_1), .n2376(n2376), .ram_s_186_0(ram_s_186_0), 
            .n2375(n2375), .ram_s_185_7(ram_s_185_7), .n2374(n2374), .ram_s_185_6(ram_s_185_6), 
            .n2373(n2373), .ram_s_185_5(ram_s_185_5), .n2372(n2372), .ram_s_185_4(ram_s_185_4), 
            .n2371(n2371), .n2370(n2370), .ram_s_185_2(ram_s_185_2), .n2369(n2369), 
            .ram_s_185_1(ram_s_185_1), .n2368(n2368), .ram_s_185_0(ram_s_185_0), 
            .n2295(n2295), .ram_s_175_7(ram_s_175_7), .n2294(n2294), .ram_s_175_6(ram_s_175_6), 
            .n2293(n2293), .ram_s_175_5(ram_s_175_5), .n2292(n2292), .ram_s_175_4(ram_s_175_4), 
            .n2291(n2291), .ram_s_175_3(ram_s_175_3), .n2290(n2290), .ram_s_175_2(ram_s_175_2), 
            .n2289(n2289), .ram_s_175_1(ram_s_175_1), .n2288(n2288), .ram_s_175_0(ram_s_175_0), 
            .n2279(n2279), .ram_s_173_7(ram_s_173_7), .n2278(n2278), .ram_s_173_6(ram_s_173_6), 
            .n2277(n2277), .ram_s_173_5(ram_s_173_5), .n2276(n2276), .ram_s_173_4(ram_s_173_4), 
            .n2275(n2275), .ram_s_173_3(ram_s_173_3), .n2274(n2274), .ram_s_173_2(ram_s_173_2), 
            .n2273(n2273), .ram_s_173_1(ram_s_173_1), .n2272(n2272), .ram_s_173_0(ram_s_173_0), 
            .n2271(n2271), .ram_s_172_7(ram_s_172_7), .n2270(n2270), .ram_s_172_6(ram_s_172_6), 
            .n2269(n2269), .ram_s_172_5(ram_s_172_5), .n2268(n2268), .ram_s_172_4(ram_s_172_4), 
            .n2267(n2267), .ram_s_172_3(ram_s_172_3), .n2266(n2266), .ram_s_172_2(ram_s_172_2), 
            .n2265(n2265), .ram_s_172_1(ram_s_172_1), .n2264(n2264), .ram_s_172_0(ram_s_172_0), 
            .n2263(n2263), .ram_s_171_7(ram_s_171_7), .n2262(n2262), .ram_s_171_6(ram_s_171_6), 
            .n2261(n2261), .n2260(n2260), .ram_s_171_4(ram_s_171_4), .n2259(n2259), 
            .ram_s_171_3(ram_s_171_3), .n2258(n2258), .ram_s_171_2(ram_s_171_2), 
            .n2257(n2257), .ram_s_171_1(ram_s_171_1), .n2256(n2256), .ram_s_171_0(ram_s_171_0), 
            .n2239(n2239), .ram_s_168_7(ram_s_168_7), .n2238(n2238), .ram_s_168_6(ram_s_168_6), 
            .n2237(n2237), .n2236(n2236), .ram_s_168_4(ram_s_168_4), .n2235(n2235), 
            .ram_s_168_3(ram_s_168_3), .n2234(n2234), .ram_s_168_2(ram_s_168_2), 
            .n2233(n2233), .ram_s_168_1(ram_s_168_1), .n2232(n2232), .ram_s_168_0(ram_s_168_0), 
            .n2231(n2231), .ram_s_167_7(ram_s_167_7), .n2230(n2230), .ram_s_167_6(ram_s_167_6), 
            .n2229(n2229), .ram_s_167_5(ram_s_167_5), .n2228(n2228), .ram_s_167_4(ram_s_167_4), 
            .n2227(n2227), .ram_s_167_3(ram_s_167_3), .n2226(n2226), .ram_s_167_2(ram_s_167_2), 
            .n2225(n2225), .ram_s_167_1(ram_s_167_1), .n2224(n2224), .ram_s_167_0(ram_s_167_0), 
            .n2223(n2223), .ram_s_166_7(ram_s_166_7), .n2222(n2222), .ram_s_166_6(ram_s_166_6), 
            .n2221(n2221), .ram_s_166_5(ram_s_166_5), .n2220(n2220), .ram_s_166_4(ram_s_166_4), 
            .n2219(n2219), .ram_s_166_3(ram_s_166_3), .n2218(n2218), .ram_s_166_2(ram_s_166_2), 
            .n2217(n2217), .ram_s_166_1(ram_s_166_1), .n2216(n2216), .ram_s_166_0(ram_s_166_0), 
            .n2215(n2215), .ram_s_165_7(ram_s_165_7), .n2214(n2214), .ram_s_165_6(ram_s_165_6), 
            .n2213(n2213), .ram_s_165_5(ram_s_165_5), .n2212(n2212), .ram_s_165_4(ram_s_165_4), 
            .n2211(n2211), .ram_s_165_3(ram_s_165_3), .n2210(n2210), .ram_s_165_2(ram_s_165_2), 
            .n2209(n2209), .ram_s_165_1(ram_s_165_1), .n2208(n2208), .ram_s_165_0(ram_s_165_0), 
            .n2207(n2207), .ram_s_164_7(ram_s_164_7), .n2206(n2206), .ram_s_164_6(ram_s_164_6), 
            .n2205(n2205), .ram_s_164_5(ram_s_164_5), .n2204(n2204), .ram_s_164_4(ram_s_164_4), 
            .n2203(n2203), .ram_s_164_3(ram_s_164_3), .n2202(n2202), .ram_s_164_2(ram_s_164_2), 
            .n2201(n2201), .ram_s_164_1(ram_s_164_1), .n2200(n2200), .ram_s_164_0(ram_s_164_0), 
            .n2199(n2199), .ram_s_163_7(ram_s_163_7), .n2198(n2198), .ram_s_163_6(ram_s_163_6), 
            .n2197(n2197), .ram_s_163_5(ram_s_163_5), .n2196(n2196), .ram_s_163_4(ram_s_163_4), 
            .n2195(n2195), .ram_s_163_3(ram_s_163_3), .n2194(n2194), .ram_s_163_2(ram_s_163_2), 
            .n2193(n2193), .ram_s_163_1(ram_s_163_1), .n2192(n2192), .ram_s_163_0(ram_s_163_0), 
            .n2191(n2191), .ram_s_162_7(ram_s_162_7), .n2190(n2190), .ram_s_162_6(ram_s_162_6), 
            .n2189(n2189), .ram_s_162_5(ram_s_162_5), .n2188(n2188), .ram_s_162_4(ram_s_162_4), 
            .n2187(n2187), .ram_s_162_3(ram_s_162_3), .n2186(n2186), .ram_s_162_2(ram_s_162_2), 
            .n2185(n2185), .ram_s_162_1(ram_s_162_1), .n2184(n2184), .ram_s_162_0(ram_s_162_0), 
            .n2183(n2183), .ram_s_161_7(ram_s_161_7), .n2182(n2182), .ram_s_161_6(ram_s_161_6), 
            .n2181(n2181), .ram_s_161_5(ram_s_161_5), .n2180(n2180), .ram_s_161_4(ram_s_161_4), 
            .n2179(n2179), .ram_s_161_3(ram_s_161_3), .n2178(n2178), .ram_s_161_2(ram_s_161_2), 
            .n2177(n2177), .ram_s_161_1(ram_s_161_1), .n2176(n2176), .ram_s_161_0(ram_s_161_0), 
            .n2175(n2175), .ram_s_160_7(ram_s_160_7), .n2174(n2174), .ram_s_160_6(ram_s_160_6), 
            .n2173(n2173), .ram_s_160_5(ram_s_160_5), .n2172(n2172), .ram_s_160_4(ram_s_160_4), 
            .n2171(n2171), .ram_s_160_3(ram_s_160_3), .n2170(n2170), .ram_s_160_2(ram_s_160_2), 
            .n2169(n2169), .ram_s_160_1(ram_s_160_1), .n2168(n2168), .ram_s_160_0(ram_s_160_0), 
            .n2031(n2031), .n2030(n2030), .ram_s_142_6(ram_s_142_6), .n2029(n2029), 
            .n2028(n2028), .ram_s_142_4(ram_s_142_4), .n2027(n2027), .n2026(n2026), 
            .ram_s_142_2(ram_s_142_2), .n2025(n2025), .ram_s_142_1(ram_s_142_1), 
            .n2024(n2024), .ram_s_142_0(ram_s_142_0), .n2023(n2023), .n2022(n2022), 
            .ram_s_141_6(ram_s_141_6), .n2021(n2021), .n2020(n2020), .ram_s_141_4(ram_s_141_4), 
            .n2019(n2019), .n2018(n2018), .ram_s_141_2(ram_s_141_2), .n2017(n2017), 
            .ram_s_141_1(ram_s_141_1), .n2016(n2016), .ram_s_141_0(ram_s_141_0), 
            .n2015(n2015), .n2014(n2014), .ram_s_140_6(ram_s_140_6), .n2013(n2013), 
            .n2012(n2012), .ram_s_140_4(ram_s_140_4), .n2011(n2011), .n2010(n2010), 
            .ram_s_140_2(ram_s_140_2), .n2009(n2009), .ram_s_140_1(ram_s_140_1), 
            .n2008(n2008), .ram_s_140_0(ram_s_140_0), .n2007(n2007), .ram_s_139_7(ram_s_139_7), 
            .n2006(n2006), .ram_s_139_6(ram_s_139_6), .n2005(n2005), .ram_s_139_5(ram_s_139_5), 
            .n2004(n2004), .ram_s_139_4(ram_s_139_4), .n2003(n2003), .ram_s_139_3(ram_s_139_3), 
            .n2002(n2002), .ram_s_139_2(ram_s_139_2), .n2001(n2001), .n2000(n2000), 
            .n1983(n1983), .ram_s_136_7(ram_s_136_7), .n1982(n1982), .ram_s_136_6(ram_s_136_6), 
            .n1981(n1981), .ram_s_136_5(ram_s_136_5), .n1980(n1980), .ram_s_136_4(ram_s_136_4), 
            .n1979(n1979), .ram_s_136_3(ram_s_136_3), .n1978(n1978), .ram_s_136_2(ram_s_136_2), 
            .n1977(n1977), .n1976(n1976), .n1975(n1975), .ram_s_135_7(ram_s_135_7), 
            .n1974(n1974), .ram_s_135_6(ram_s_135_6), .n1973(n1973), .n1972(n1972), 
            .ram_s_135_4(ram_s_135_4), .n1971(n1971), .ram_s_135_3(ram_s_135_3), 
            .n1970(n1970), .ram_s_135_2(ram_s_135_2), .n1969(n1969), .ram_s_135_1(ram_s_135_1), 
            .n1968(n1968), .n1967(n1967), .ram_s_134_7(ram_s_134_7), .n1966(n1966), 
            .ram_s_134_6(ram_s_134_6), .n1965(n1965), .n1964(n1964), .ram_s_134_4(ram_s_134_4), 
            .n1963(n1963), .ram_s_134_3(ram_s_134_3), .n1962(n1962), .ram_s_134_2(ram_s_134_2), 
            .n1961(n1961), .ram_s_134_1(ram_s_134_1), .n1960(n1960), .n1959(n1959), 
            .ram_s_133_7(ram_s_133_7), .n1958(n1958), .ram_s_133_6(ram_s_133_6), 
            .n1957(n1957), .n1956(n1956), .ram_s_133_4(ram_s_133_4), .n1955(n1955), 
            .ram_s_133_3(ram_s_133_3), .n1954(n1954), .ram_s_133_2(ram_s_133_2), 
            .n1953(n1953), .ram_s_133_1(ram_s_133_1), .n1952(n1952), .n1951(n1951), 
            .ram_s_132_7(ram_s_132_7), .n1950(n1950), .ram_s_132_6(ram_s_132_6), 
            .n1949(n1949), .n1948(n1948), .ram_s_132_4(ram_s_132_4), .n1947(n1947), 
            .ram_s_132_3(ram_s_132_3), .n1946(n1946), .ram_s_132_2(ram_s_132_2), 
            .n1945(n1945), .ram_s_132_1(ram_s_132_1), .n1944(n1944), .n1943(n1943), 
            .n1942(n1942), .ram_s_131_6(ram_s_131_6), .n1941(n1941), .ram_s_131_5(ram_s_131_5), 
            .n1940(n1940), .ram_s_131_4(ram_s_131_4), .n1939(n1939), .ram_s_131_3(ram_s_131_3), 
            .n1938(n1938), .ram_s_131_2(ram_s_131_2), .n1937(n1937), .ram_s_131_1(ram_s_131_1), 
            .n1936(n1936), .n1935(n1935), .n1934(n1934), .ram_s_130_6(ram_s_130_6), 
            .n1933(n1933), .ram_s_130_5(ram_s_130_5), .n1932(n1932), .ram_s_130_4(ram_s_130_4), 
            .n1931(n1931), .ram_s_130_3(ram_s_130_3), .n1930(n1930), .ram_s_130_2(ram_s_130_2), 
            .n1929(n1929), .ram_s_130_1(ram_s_130_1), .n1928(n1928), .n1927(n1927), 
            .n1926(n1926), .ram_s_129_6(ram_s_129_6), .n1925(n1925), .ram_s_129_5(ram_s_129_5), 
            .n1924(n1924), .ram_s_129_4(ram_s_129_4), .n1923(n1923), .ram_s_129_3(ram_s_129_3), 
            .n1922(n1922), .ram_s_129_2(ram_s_129_2), .n1921(n1921), .ram_s_129_1(ram_s_129_1), 
            .n1920(n1920), .n1919(n1919), .n1918(n1918), .ram_s_128_6(ram_s_128_6), 
            .n1917(n1917), .ram_s_128_5(ram_s_128_5), .n1916(n1916), .ram_s_128_4(ram_s_128_4), 
            .n1915(n1915), .ram_s_128_3(ram_s_128_3), .n1914(n1914), .ram_s_128_2(ram_s_128_2), 
            .n1913(n1913), .ram_s_128_1(ram_s_128_1), .n1912(n1912), .n1543(n1543), 
            .ram_s_81_7(ram_s_81_7), .n1542(n1542), .ram_s_81_6(ram_s_81_6), 
            .n1541(n1541), .n1540(n1540), .ram_s_81_4(ram_s_81_4), .n1539(n1539), 
            .ram_s_81_3(ram_s_81_3), .n1538(n1538), .ram_s_81_2(ram_s_81_2), 
            .n1537(n1537), .ram_s_81_1(ram_s_81_1), .n1536(n1536), .ram_s_81_0(ram_s_81_0), 
            .n1495(n1495), .n1494(n1494), .ram_s_75_6(ram_s_75_6), .n1493(n1493), 
            .ram_s_75_5(ram_s_75_5), .n1492(n1492), .n1491(n1491), .ram_s_75_3(ram_s_75_3), 
            .n1490(n1490), .n1489(n1489), .ram_s_75_1(ram_s_75_1), .n1488(n1488), 
            .ram_s_75_0(ram_s_75_0), .n1487(n1487), .n1486(n1486), .ram_s_74_6(ram_s_74_6), 
            .n1485(n1485), .ram_s_74_5(ram_s_74_5), .n1484(n1484), .n1483(n1483), 
            .ram_s_74_3(ram_s_74_3), .n1482(n1482), .n1481(n1481), .ram_s_74_1(ram_s_74_1), 
            .n1480(n1480), .ram_s_74_0(ram_s_74_0), .n1479(n1479), .n1478(n1478), 
            .ram_s_73_6(ram_s_73_6), .n1477(n1477), .ram_s_73_5(ram_s_73_5), 
            .n1476(n1476), .n1475(n1475), .ram_s_73_3(ram_s_73_3), .n1474(n1474), 
            .n1473(n1473), .ram_s_73_1(ram_s_73_1), .n1472(n1472), .ram_s_73_0(ram_s_73_0), 
            .n1471(n1471), .n1470(n1470), .ram_s_72_6(ram_s_72_6), .n1469(n1469), 
            .ram_s_72_5(ram_s_72_5), .n1468(n1468), .n1467(n1467), .ram_s_72_3(ram_s_72_3), 
            .n1466(n1466), .n1465(n1465), .ram_s_72_1(ram_s_72_1), .n1464(n1464), 
            .ram_s_72_0(ram_s_72_0), .n1463(n1463), .ram_s_71_7(ram_s_71_7), 
            .n1462(n1462), .ram_s_71_6(ram_s_71_6), .n1461(n1461), .ram_s_71_5(ram_s_71_5), 
            .n1460(n1460), .n1459(n1459), .n1458(n1458), .ram_s_71_2(ram_s_71_2), 
            .n1457(n1457), .ram_s_71_1(ram_s_71_1), .n1456(n1456), .ram_s_71_0(ram_s_71_0), 
            .n1455(n1455), .ram_s_70_7(ram_s_70_7), .n1454(n1454), .ram_s_70_6(ram_s_70_6), 
            .n1453(n1453), .ram_s_70_5(ram_s_70_5), .n1452(n1452), .n1451(n1451), 
            .n1450(n1450), .ram_s_70_2(ram_s_70_2), .n1449(n1449), .ram_s_70_1(ram_s_70_1), 
            .n1448(n1448), .ram_s_70_0(ram_s_70_0), .n1447(n1447), .ram_s_69_7(ram_s_69_7), 
            .n1446(n1446), .ram_s_69_6(ram_s_69_6), .n1445(n1445), .ram_s_69_5(ram_s_69_5), 
            .n1444(n1444), .n1443(n1443), .n1442(n1442), .ram_s_69_2(ram_s_69_2), 
            .n1441(n1441), .ram_s_69_1(ram_s_69_1), .n1440(n1440), .ram_s_69_0(ram_s_69_0), 
            .n1439(n1439), .ram_s_68_7(ram_s_68_7), .n1438(n1438), .ram_s_68_6(ram_s_68_6), 
            .n1437(n1437), .ram_s_68_5(ram_s_68_5), .n1436(n1436), .n1435(n1435), 
            .n1434(n1434), .ram_s_68_2(ram_s_68_2), .n1433(n1433), .ram_s_68_1(ram_s_68_1), 
            .n1432(n1432), .ram_s_68_0(ram_s_68_0), .n1431(n1431), .ram_s_67_7(ram_s_67_7), 
            .n1430(n1430), .ram_s_67_6(ram_s_67_6), .n1429(n1429), .ram_s_67_5(ram_s_67_5), 
            .n1428(n1428), .n1427(n1427), .ram_s_67_3(ram_s_67_3), .n1426(n1426), 
            .ram_s_67_2(ram_s_67_2), .n1425(n1425), .ram_s_67_1(ram_s_67_1), 
            .n1424(n1424), .n1423(n1423), .ram_s_66_7(ram_s_66_7), .n1422(n1422), 
            .ram_s_66_6(ram_s_66_6), .n1421(n1421), .ram_s_66_5(ram_s_66_5), 
            .n1420(n1420), .n1419(n1419), .ram_s_66_3(ram_s_66_3), .n1418(n1418), 
            .ram_s_66_2(ram_s_66_2), .n1417(n1417), .ram_s_66_1(ram_s_66_1), 
            .n1416(n1416), .n1415(n1415), .ram_s_65_7(ram_s_65_7), .n1414(n1414), 
            .ram_s_65_6(ram_s_65_6), .n1413(n1413), .ram_s_65_5(ram_s_65_5), 
            .n1412(n1412), .n1411(n1411), .ram_s_65_3(ram_s_65_3), .n1410(n1410), 
            .ram_s_65_2(ram_s_65_2), .n1409(n1409), .ram_s_65_1(ram_s_65_1), 
            .n1408(n1408), .n1407(n1407), .ram_s_64_7(ram_s_64_7), .n1406(n1406), 
            .ram_s_64_6(ram_s_64_6), .n1405(n1405), .ram_s_64_5(ram_s_64_5), 
            .n1404(n1404), .n1403(n1403), .ram_s_64_3(ram_s_64_3), .n1402(n1402), 
            .ram_s_64_2(ram_s_64_2), .n1401(n1401), .ram_s_64_1(ram_s_64_1), 
            .n1400(n1400), .n1399(n1399), .ram_s_63_7(ram_s_63_7), .n1398(n1398), 
            .ram_s_63_6(ram_s_63_6), .n1397(n1397), .ram_s_63_5(ram_s_63_5), 
            .n1396(n1396), .n1395(n1395), .ram_s_63_3(ram_s_63_3), .n1394(n1394), 
            .ram_s_63_2(ram_s_63_2), .n1393(n1393), .ram_s_63_1(ram_s_63_1), 
            .n1392(n1392), .n1391(n1391), .ram_s_62_7(ram_s_62_7), .n1390(n1390), 
            .ram_s_62_6(ram_s_62_6), .n1389(n1389), .ram_s_62_5(ram_s_62_5), 
            .n1388(n1388), .n1387(n1387), .ram_s_62_3(ram_s_62_3), .n1386(n1386), 
            .ram_s_62_2(ram_s_62_2), .n1385(n1385), .ram_s_62_1(ram_s_62_1), 
            .n1384(n1384), .n1359(n1359), .ram_s_58_7(ram_s_58_7), .n1358(n1358), 
            .ram_s_58_6(ram_s_58_6), .n1357(n1357), .n1356(n1356), .ram_s_58_4(ram_s_58_4), 
            .n1355(n1355), .ram_s_58_3(ram_s_58_3), .n1354(n1354), .ram_s_58_2(ram_s_58_2), 
            .n1353(n1353), .ram_s_58_1(ram_s_58_1), .n1352(n1352), .n1351(n1351), 
            .ram_s_57_7(ram_s_57_7), .n1350(n1350), .ram_s_57_6(ram_s_57_6), 
            .n1349(n1349), .n1348(n1348), .ram_s_57_4(ram_s_57_4), .n1347(n1347), 
            .ram_s_57_3(ram_s_57_3), .n1346(n1346), .ram_s_57_2(ram_s_57_2), 
            .n1345(n1345), .ram_s_57_1(ram_s_57_1), .n1344(n1344), .n1271(n1271), 
            .ram_s_47_7(ram_s_47_7), .n1270(n1270), .ram_s_47_6(ram_s_47_6), 
            .n1269(n1269), .ram_s_47_5(ram_s_47_5), .n1268(n1268), .ram_s_47_4(ram_s_47_4), 
            .n1267(n1267), .ram_s_47_3(ram_s_47_3), .n1266(n1266), .n1265(n1265), 
            .ram_s_47_1(ram_s_47_1), .n1264(n1264), .ram_s_47_0(ram_s_47_0), 
            .n1255(n1255), .ram_s_45_7(ram_s_45_7), .n1254(n1254), .ram_s_45_6(ram_s_45_6), 
            .n1253(n1253), .ram_s_45_5(ram_s_45_5), .n1252(n1252), .ram_s_45_4(ram_s_45_4), 
            .n1251(n1251), .ram_s_45_3(ram_s_45_3), .n1250(n1250), .n1249(n1249), 
            .ram_s_45_1(ram_s_45_1), .n1248(n1248), .ram_s_45_0(ram_s_45_0), 
            .n1247(n1247), .ram_s_44_7(ram_s_44_7), .n1246(n1246), .ram_s_44_6(ram_s_44_6), 
            .n1245(n1245), .ram_s_44_5(ram_s_44_5), .n1244(n1244), .ram_s_44_4(ram_s_44_4), 
            .n1243(n1243), .ram_s_44_3(ram_s_44_3), .n1242(n1242), .n1241(n1241), 
            .ram_s_44_1(ram_s_44_1), .n1240(n1240), .ram_s_44_0(ram_s_44_0), 
            .n1239(n1239), .n1238(n1238), .ram_s_43_6(ram_s_43_6), .n1237(n1237), 
            .ram_s_43_5(ram_s_43_5), .n1236(n1236), .ram_s_43_4(ram_s_43_4), 
            .n1235(n1235), .ram_s_43_3(ram_s_43_3), .n1234(n1234), .n1233(n1233), 
            .n1232(n1232), .ram_s_43_0(ram_s_43_0), .n1215(n1215), .n1214(n1214), 
            .ram_s_40_6(ram_s_40_6), .n1213(n1213), .ram_s_40_5(ram_s_40_5), 
            .n1212(n1212), .ram_s_40_4(ram_s_40_4), .n1211(n1211), .ram_s_40_3(ram_s_40_3), 
            .n1210(n1210), .n1209(n1209), .n1208(n1208), .ram_s_40_0(ram_s_40_0), 
            .n1207(n1207), .n1206(n1206), .ram_s_39_6(ram_s_39_6), .n1205(n1205), 
            .ram_s_39_5(ram_s_39_5), .n1204(n1204), .ram_s_39_4(ram_s_39_4), 
            .n1203(n1203), .ram_s_39_3(ram_s_39_3), .n1202(n1202), .ram_s_39_2(ram_s_39_2), 
            .n1201(n1201), .ram_s_39_1(ram_s_39_1), .n1200(n1200), .n1199(n1199), 
            .n1198(n1198), .ram_s_38_6(ram_s_38_6), .n1197(n1197), .ram_s_38_5(ram_s_38_5), 
            .n1196(n1196), .ram_s_38_4(ram_s_38_4), .n1195(n1195), .ram_s_38_3(ram_s_38_3), 
            .n1194(n1194), .ram_s_38_2(ram_s_38_2), .n1193(n1193), .ram_s_38_1(ram_s_38_1), 
            .n1192(n1192), .n1191(n1191), .n1190(n1190), .ram_s_37_6(ram_s_37_6), 
            .n1189(n1189), .ram_s_37_5(ram_s_37_5), .n1188(n1188), .ram_s_37_4(ram_s_37_4), 
            .n1187(n1187), .ram_s_37_3(ram_s_37_3), .n1186(n1186), .ram_s_37_2(ram_s_37_2), 
            .n1185(n1185), .ram_s_37_1(ram_s_37_1), .n1184(n1184), .n1183(n1183), 
            .n1182(n1182), .ram_s_36_6(ram_s_36_6), .n1181(n1181), .ram_s_36_5(ram_s_36_5), 
            .n1180(n1180), .ram_s_36_4(ram_s_36_4), .n1179(n1179), .ram_s_36_3(ram_s_36_3), 
            .n1178(n1178), .ram_s_36_2(ram_s_36_2), .n1177(n1177), .ram_s_36_1(ram_s_36_1), 
            .n1176(n1176), .n1175(n1175), .n1174(n1174), .ram_s_35_6(ram_s_35_6), 
            .n1173(n1173), .ram_s_35_5(ram_s_35_5), .n1172(n1172), .ram_s_35_4(ram_s_35_4), 
            .n1171(n1171), .ram_s_35_3(ram_s_35_3), .n1170(n1170), .n1169(n1169), 
            .n1168(n1168), .ram_s_35_0(ram_s_35_0), .n1167(n1167), .n1166(n1166), 
            .ram_s_34_6(ram_s_34_6), .n1165(n1165), .ram_s_34_5(ram_s_34_5), 
            .n1164(n1164), .ram_s_34_4(ram_s_34_4), .n1163(n1163), .ram_s_34_3(ram_s_34_3), 
            .n1162(n1162), .n1161(n1161), .n1160(n1160), .ram_s_34_0(ram_s_34_0), 
            .n1159(n1159), .n1158(n1158), .ram_s_33_6(ram_s_33_6), .n1157(n1157), 
            .ram_s_33_5(ram_s_33_5), .n1156(n1156), .ram_s_33_4(ram_s_33_4), 
            .n1155(n1155), .ram_s_33_3(ram_s_33_3), .n1154(n1154), .n1153(n1153), 
            .n1152(n1152), .ram_s_33_0(ram_s_33_0), .n1151(n1151), .n1150(n1150), 
            .ram_s_32_6(ram_s_32_6), .n1149(n1149), .ram_s_32_5(ram_s_32_5), 
            .n1148(n1148), .ram_s_32_4(ram_s_32_4), .n1147(n1147), .ram_s_32_3(ram_s_32_3), 
            .n1146(n1146), .n1145(n1145), .n1144(n1144), .ram_s_32_0(ram_s_32_0), 
            .n1051(n1051), .n1047(n1047), .n1046(n1046), .n1045(n1045), 
            .ram_s_0_2(ram_s_0_2), .n1044(n1044), .ram_s_12_3(ram_s_12_3), 
            .n1043(n1043), .n1042(n1042), .ram_s_11_1(ram_s_11_1), .n1041(n1041), 
            .n1040(n1040), .ram_s_12_1(ram_s_12_1), .n1038(n1038), .ram_s_11_4(ram_s_11_4), 
            .n182(n182), .n1037(n1037), .ram_s_12_4(ram_s_12_4), .n54(n54), 
            .n1036(n1036), .ram_s_11_7(ram_s_11_7), .n183(n183), .n1035(n1035), 
            .n55(n55), .n1034(n1034), .ram_s_12_7(ram_s_12_7), .n184(n184), 
            .n1033(n1033), .ram_s_12_2(ram_s_12_2), .n56(n56), .n1032(n1032), 
            .ram_s_11_5(ram_s_11_5), .n185(n185), .n1031(n1031), .n57(n57), 
            .n1030(n1030), .ram_s_12_0(ram_s_12_0), .n186(n186), .n1029(n1029), 
            .ram_s_11_3(ram_s_11_3), .n58(n58), .n187(n187), .n59(n59), 
            .n188(n188), .n60(n60), .n189(n189), .n61(n61), .n190(n190), 
            .n62(n62), .n191(n191), .n63(n63), .n192(n192), .n1017(n1017), 
            .ram_s_0_3(ram_s_0_3), .n64(n64), .n1016(n1016), .ram_s_0_4(ram_s_0_4), 
            .n193(n193), .n1015(n1015), .ram_s_0_5(ram_s_0_5), .n65(n65), 
            .n1014(n1014), .ram_s_0_6(ram_s_0_6), .n194(n194), .n1013(n1013), 
            .n66(n66), .n1012(n1012), .n195(n195), .n1011(n1011), .n67(n67), 
            .n1010(n1010), .ram_s_1_2(ram_s_1_2), .n1009(n1009), .ram_s_1_3(ram_s_1_3), 
            .n1008(n1008), .ram_s_1_4(ram_s_1_4), .n1007(n1007), .ram_s_1_5(ram_s_1_5), 
            .n1006(n1006), .ram_s_4_4(ram_s_4_4), .n1005(n1005), .n1004(n1004), 
            .n1003(n1003), .ram_s_5_0(ram_s_5_0), .n1002(n1002), .ram_s_4_6(ram_s_4_6), 
            .n1001(n1001), .ram_s_5_1(ram_s_5_1), .n998(n998), .ram_s_8_5(ram_s_8_5), 
            .n997(n997), .n996(n996), .n995(n995), .ram_s_7_4(ram_s_7_4), 
            .n994(n994), .ram_s_7_1(ram_s_7_1), .n993(n993), .ram_s_6_6(ram_s_6_6), 
            .n992(n992), .ram_s_6_3(ram_s_6_3), .n989(n989), .n988(n988), 
            .ram_s_8_3(ram_s_8_3), .n987(n987), .ram_s_8_0(ram_s_8_0), 
            .n986(n986), .n199(n199), .n985(n985), .ram_s_7_2(ram_s_7_2), 
            .n71(n71), .n984(n984), .n200(n200), .n983(n983), .ram_s_6_4(ram_s_6_4), 
            .n72(n72), .n980(n980), .ram_s_8_7(ram_s_8_7), .n979(n979), 
            .ram_s_8_4(ram_s_8_4), .n978(n978), .ram_s_8_1(ram_s_8_1), 
            .n977(n977), .ram_s_7_6(ram_s_7_6), .n976(n976), .ram_s_7_3(ram_s_7_3), 
            .n975(n975), .ram_s_7_0(ram_s_7_0), .n974(n974), .n973(n973), 
            .ram_s_1_6(ram_s_1_6), .n972(n972), .n971(n971), .n970(n970), 
            .n969(n969), .ram_s_2_2(ram_s_2_2), .n968(n968), .ram_s_2_3(ram_s_2_3), 
            .n967(n967), .ram_s_2_4(ram_s_2_4), .n966(n966), .ram_s_2_5(ram_s_2_5), 
            .n965(n965), .ram_s_2_6(ram_s_2_6), .n964(n964), .n963(n963), 
            .n962(n962), .n961(n961), .ram_s_3_2(ram_s_3_2), .n960(n960), 
            .ram_s_3_3(ram_s_3_3), .n959(n959), .ram_s_3_4(ram_s_3_4), 
            .n958(n958), .ram_s_3_5(ram_s_3_5), .n957(n957), .ram_s_14_7(ram_s_14_7), 
            .n952(n952), .ram_s_3_6(ram_s_3_6), .n950(n950), .n946(n946), 
            .ram_s_4_0(ram_s_4_0), .n944(n944), .ram_s_4_1(ram_s_4_1), 
            .n941(n941), .ram_s_4_2(ram_s_4_2), .n940(n940), .ram_s_5_2(ram_s_5_2), 
            .n939(n939), .ram_s_5_3(ram_s_5_3), .n935(n935), .n934(n934), 
            .ram_s_6_0(ram_s_6_0), .n933(n933), .ram_s_6_1(ram_s_6_1), 
            .n932(n932), .ram_s_6_2(ram_s_6_2), .n931(n931), .ram_s_5_6(ram_s_5_6), 
            .n930(n930), .n927(n927), .ram_s_4_3(ram_s_4_3), .n926(n926), 
            .n925(n925), .ram_s_13_3(ram_s_13_3), .n924(n924), .ram_s_13_4(ram_s_13_4), 
            .n923(n923), .n210(n210), .n82(n82), .n212(n212), .n84(n84), 
            .n213(n213), .n85(n85), .n214(n214), .n86(n86), .n217(n217), 
            .n89(n89), .n218(n218), .n90(n90), .n219(n219), .n91(n91), 
            .n220(n220), .n92(n92), .n221(n221), .n93(n93), .n222(n222), 
            .n94(n94), .n223(n223), .n95(n95), .n224(n224), .n96(n96), 
            .n225(n225), .n97(n97), .n918(n918), .ram_s_13_7(ram_s_13_7), 
            .n917(n917), .ram_s_14_0(ram_s_14_0), .n916(n916), .ram_s_14_1(ram_s_14_1), 
            .spm_enable(spm_enable), .n244(n244), .n116(n116), .n115(n115), 
            .n243(n243), .n245(n245), .n117(n117), .n246(n246), .n118(n118), 
            .n48(n48), .n176(n176), .n249(n249), .n121(n121), .n250(n250), 
            .n122(n122), .n251(n251), .n123(n123), .n252(n252), .n124(n124), 
            .n253(n253), .n125(n125), .n254(n254), .n126(n126), .n255(n255), 
            .n127(n127), .n256(n256), .n128(n128), .n257(n257), .n129(n129), 
            .ram_s_14_2(ram_s_14_2), .ram_s_13_2(ram_s_13_2), .ram_s_11_0(ram_s_11_0), 
            .n911(n911), .n909(n909), .n908(n908), .ram_s_14_3(ram_s_14_3), 
            .n907(n907), .ram_s_13_1(ram_s_13_1), .n906(n906), .n904(n904), 
            .ram_s_13_0(ram_s_13_0), .n901(n901), .ram_s_5_4(ram_s_5_4), 
            .n899(n899));   // src/spm_with_output_reg.vhd(145[12:15])
    
endmodule
//
// Verilog Description of module \ram(8,8) 
//

module \ram(8,8)  (port_id, ram_s_70_3, ram_s_71_3, ram_s_69_3, ram_s_68_3, 
            \sx[7] , \sx[6] , \sx[5] , \sx[4] , \register_vector[10] , 
            ram_s_34_7, ram_s_35_7, ram_s_33_7, ram_s_32_7, \register_vector[9] , 
            ram_s_11_6, ram_s_8_6, \register_vector[11] , ram_s_62_4, 
            ram_s_63_4, ram_s_2_7, ram_s_3_7, ram_s_1_7, ram_s_0_7, 
            ram_s_66_4, ram_s_67_4, ram_s_65_4, ram_s_64_4, \register_vector[8] , 
            ram_s_142_3, ram_s_141_3, ram_s_140_3, CLK_3P3_MHZ_c, ram_s_209_3, 
            ram_s_130_0, ram_s_131_0, ram_s_129_0, ram_s_128_0, ram_s_70_4, 
            ram_s_71_4, ram_s_69_4, ram_s_68_4, ram_s_171_5, ram_s_168_5, 
            ram_s_14_6, ram_s_13_6, ram_s_12_6, ram_s_202_1, ram_s_203_1, 
            ram_s_6_5, ram_s_7_5, ram_s_14_5, ram_s_5_5, ram_s_4_5, 
            ram_s_13_5, ram_s_12_5, ram_s_43_2, ram_s_2_0, ram_s_3_0, 
            ram_s_2_1, ram_s_3_1, ram_s_1_0, ram_s_0_0, ram_s_66_0, 
            ram_s_67_0, ram_s_34_1, ram_s_35_1, ram_s_33_1, ram_s_32_1, 
            ram_s_201_1, ram_s_200_1, ram_s_1_1, ram_s_0_1, ram_s_65_0, 
            ram_s_64_0, ram_s_11_2, ram_s_8_2, ram_s_38_0, ram_s_39_0, 
            ram_s_40_2, ram_s_74_7, ram_s_75_7, ram_s_73_7, ram_s_72_7, 
            ram_s_130_7, ram_s_131_7, ram_s_129_7, ram_s_128_7, ram_s_37_0, 
            ram_s_36_0, ram_s_142_5, ram_s_141_5, ram_s_140_5, ram_s_62_0, 
            ram_s_63_0, ram_s_194_1, ram_s_195_1, ram_s_193_1, ram_s_192_1, 
            ram_s_74_4, ram_s_75_4, ram_s_73_4, ram_s_72_4, ram_s_43_7, 
            ram_s_40_7, ram_s_74_2, ram_s_75_2, ram_s_73_2, ram_s_72_2, 
            ram_s_186_3, ram_s_185_3, ram_s_190_2, ram_s_191_2, ram_s_43_1, 
            wea, ram_s_40_1, ram_s_6_7, ram_s_7_7, ram_s_134_0, ram_s_135_0, 
            ram_s_5_7, ram_s_4_7, ram_s_133_0, ram_s_132_0, ram_s_34_2, 
            ram_s_35_2, ram_s_58_5, ram_s_58_0, ram_s_57_0, ram_s_139_0, 
            ram_s_136_0, ram_s_190_5, ram_s_191_5, ram_s_57_5, ram_s_33_2, 
            ram_s_32_2, ram_s_142_7, ram_s_141_7, ram_s_140_7, ram_s_81_5, 
            ram_s_190_1, ram_s_191_1, ram_s_139_1, ram_s_136_1, ram_s_38_7, 
            ram_s_39_7, ram_s_37_7, ram_s_36_7, n893, ram_s_14_4, 
            ram_s_190_7, ram_s_191_7, ram_s_47_2, spm_ram_data, ram_s_45_2, 
            ram_s_44_2, ram_s_134_5, ram_s_135_5, ram_s_133_5, ram_s_132_5, 
            n2567, ram_s_209_7, n2566, ram_s_209_6, n2565, ram_s_209_5, 
            n2564, ram_s_209_4, n2563, n2562, ram_s_209_2, n2561, 
            ram_s_209_1, n2560, ram_s_209_0, n2519, ram_s_203_7, n2518, 
            ram_s_203_6, n2517, ram_s_203_5, n2516, ram_s_203_4, n2515, 
            ram_s_203_3, n2514, ram_s_203_2, n2513, n2512, ram_s_203_0, 
            n2511, ram_s_202_7, n2510, ram_s_202_6, n2509, ram_s_202_5, 
            n2508, ram_s_202_4, n2507, ram_s_202_3, n2506, ram_s_202_2, 
            n2505, n2504, ram_s_202_0, n2503, ram_s_201_7, n2502, 
            ram_s_201_6, n2501, ram_s_201_5, n2500, ram_s_201_4, n2499, 
            ram_s_201_3, n2498, ram_s_201_2, n2497, n2496, ram_s_201_0, 
            n2495, ram_s_200_7, n2494, ram_s_200_6, n2493, ram_s_200_5, 
            n2492, ram_s_200_4, n2491, ram_s_200_3, n2490, ram_s_200_2, 
            n2489, n2488, ram_s_200_0, n2487, ram_s_199_7, n2486, 
            ram_s_199_6, n2485, ram_s_199_5, n2484, ram_s_199_4, n2483, 
            ram_s_199_3, n2482, ram_s_199_2, n2481, ram_s_199_1, n2480, 
            ram_s_199_0, n2479, ram_s_198_7, n2478, ram_s_198_6, n2477, 
            ram_s_198_5, n2476, ram_s_198_4, n2475, ram_s_198_3, n2474, 
            ram_s_198_2, n2473, ram_s_198_1, n2472, ram_s_198_0, n2471, 
            ram_s_197_7, n2470, ram_s_197_6, n2469, ram_s_197_5, n2468, 
            ram_s_197_4, n2467, ram_s_197_3, n2466, ram_s_197_2, n2465, 
            ram_s_197_1, n2464, ram_s_197_0, n2463, ram_s_196_7, n2462, 
            ram_s_196_6, n2461, ram_s_196_5, n2460, ram_s_196_4, n2459, 
            ram_s_196_3, n2458, ram_s_196_2, n2457, ram_s_196_1, n2456, 
            ram_s_196_0, n2455, ram_s_195_7, n2454, ram_s_195_6, n2453, 
            ram_s_195_5, n2452, ram_s_195_4, n2451, ram_s_195_3, n2450, 
            ram_s_195_2, n2449, n2448, ram_s_195_0, n2447, ram_s_194_7, 
            n2446, ram_s_194_6, n2445, ram_s_194_5, n2444, ram_s_194_4, 
            n2443, ram_s_194_3, n2442, ram_s_194_2, n2441, n2440, 
            ram_s_194_0, n2439, ram_s_193_7, n2438, ram_s_193_6, n2437, 
            ram_s_193_5, n2436, ram_s_193_4, n2435, ram_s_193_3, n2434, 
            ram_s_193_2, n2433, n2432, ram_s_193_0, n2431, ram_s_192_7, 
            n2430, ram_s_192_6, n2429, ram_s_192_5, n2428, ram_s_192_4, 
            n2427, ram_s_192_3, n2426, ram_s_192_2, n2425, n2424, 
            ram_s_192_0, n2423, n2422, ram_s_191_6, n2421, n2420, 
            ram_s_191_4, n2419, ram_s_191_3, n2418, n2417, n2416, 
            ram_s_191_0, n2415, n2414, ram_s_190_6, n2413, n2412, 
            ram_s_190_4, n2411, ram_s_190_3, n2410, n2409, n2408, 
            ram_s_190_0, n2383, ram_s_186_7, n2382, ram_s_186_6, n2381, 
            ram_s_186_5, n2380, ram_s_186_4, n2379, n2378, ram_s_186_2, 
            n2377, ram_s_186_1, n2376, ram_s_186_0, n2375, ram_s_185_7, 
            n2374, ram_s_185_6, n2373, ram_s_185_5, n2372, ram_s_185_4, 
            n2371, n2370, ram_s_185_2, n2369, ram_s_185_1, n2368, 
            ram_s_185_0, n2295, ram_s_175_7, n2294, ram_s_175_6, n2293, 
            ram_s_175_5, n2292, ram_s_175_4, n2291, ram_s_175_3, n2290, 
            ram_s_175_2, n2289, ram_s_175_1, n2288, ram_s_175_0, n2279, 
            ram_s_173_7, n2278, ram_s_173_6, n2277, ram_s_173_5, n2276, 
            ram_s_173_4, n2275, ram_s_173_3, n2274, ram_s_173_2, n2273, 
            ram_s_173_1, n2272, ram_s_173_0, n2271, ram_s_172_7, n2270, 
            ram_s_172_6, n2269, ram_s_172_5, n2268, ram_s_172_4, n2267, 
            ram_s_172_3, n2266, ram_s_172_2, n2265, ram_s_172_1, n2264, 
            ram_s_172_0, n2263, ram_s_171_7, n2262, ram_s_171_6, n2261, 
            n2260, ram_s_171_4, n2259, ram_s_171_3, n2258, ram_s_171_2, 
            n2257, ram_s_171_1, n2256, ram_s_171_0, n2239, ram_s_168_7, 
            n2238, ram_s_168_6, n2237, n2236, ram_s_168_4, n2235, 
            ram_s_168_3, n2234, ram_s_168_2, n2233, ram_s_168_1, n2232, 
            ram_s_168_0, n2231, ram_s_167_7, n2230, ram_s_167_6, n2229, 
            ram_s_167_5, n2228, ram_s_167_4, n2227, ram_s_167_3, n2226, 
            ram_s_167_2, n2225, ram_s_167_1, n2224, ram_s_167_0, n2223, 
            ram_s_166_7, n2222, ram_s_166_6, n2221, ram_s_166_5, n2220, 
            ram_s_166_4, n2219, ram_s_166_3, n2218, ram_s_166_2, n2217, 
            ram_s_166_1, n2216, ram_s_166_0, n2215, ram_s_165_7, n2214, 
            ram_s_165_6, n2213, ram_s_165_5, n2212, ram_s_165_4, n2211, 
            ram_s_165_3, n2210, ram_s_165_2, n2209, ram_s_165_1, n2208, 
            ram_s_165_0, n2207, ram_s_164_7, n2206, ram_s_164_6, n2205, 
            ram_s_164_5, n2204, ram_s_164_4, n2203, ram_s_164_3, n2202, 
            ram_s_164_2, n2201, ram_s_164_1, n2200, ram_s_164_0, n2199, 
            ram_s_163_7, n2198, ram_s_163_6, n2197, ram_s_163_5, n2196, 
            ram_s_163_4, n2195, ram_s_163_3, n2194, ram_s_163_2, n2193, 
            ram_s_163_1, n2192, ram_s_163_0, n2191, ram_s_162_7, n2190, 
            ram_s_162_6, n2189, ram_s_162_5, n2188, ram_s_162_4, n2187, 
            ram_s_162_3, n2186, ram_s_162_2, n2185, ram_s_162_1, n2184, 
            ram_s_162_0, n2183, ram_s_161_7, n2182, ram_s_161_6, n2181, 
            ram_s_161_5, n2180, ram_s_161_4, n2179, ram_s_161_3, n2178, 
            ram_s_161_2, n2177, ram_s_161_1, n2176, ram_s_161_0, n2175, 
            ram_s_160_7, n2174, ram_s_160_6, n2173, ram_s_160_5, n2172, 
            ram_s_160_4, n2171, ram_s_160_3, n2170, ram_s_160_2, n2169, 
            ram_s_160_1, n2168, ram_s_160_0, n2031, n2030, ram_s_142_6, 
            n2029, n2028, ram_s_142_4, n2027, n2026, ram_s_142_2, 
            n2025, ram_s_142_1, n2024, ram_s_142_0, n2023, n2022, 
            ram_s_141_6, n2021, n2020, ram_s_141_4, n2019, n2018, 
            ram_s_141_2, n2017, ram_s_141_1, n2016, ram_s_141_0, n2015, 
            n2014, ram_s_140_6, n2013, n2012, ram_s_140_4, n2011, 
            n2010, ram_s_140_2, n2009, ram_s_140_1, n2008, ram_s_140_0, 
            n2007, ram_s_139_7, n2006, ram_s_139_6, n2005, ram_s_139_5, 
            n2004, ram_s_139_4, n2003, ram_s_139_3, n2002, ram_s_139_2, 
            n2001, n2000, n1983, ram_s_136_7, n1982, ram_s_136_6, 
            n1981, ram_s_136_5, n1980, ram_s_136_4, n1979, ram_s_136_3, 
            n1978, ram_s_136_2, n1977, n1976, n1975, ram_s_135_7, 
            n1974, ram_s_135_6, n1973, n1972, ram_s_135_4, n1971, 
            ram_s_135_3, n1970, ram_s_135_2, n1969, ram_s_135_1, n1968, 
            n1967, ram_s_134_7, n1966, ram_s_134_6, n1965, n1964, 
            ram_s_134_4, n1963, ram_s_134_3, n1962, ram_s_134_2, n1961, 
            ram_s_134_1, n1960, n1959, ram_s_133_7, n1958, ram_s_133_6, 
            n1957, n1956, ram_s_133_4, n1955, ram_s_133_3, n1954, 
            ram_s_133_2, n1953, ram_s_133_1, n1952, n1951, ram_s_132_7, 
            n1950, ram_s_132_6, n1949, n1948, ram_s_132_4, n1947, 
            ram_s_132_3, n1946, ram_s_132_2, n1945, ram_s_132_1, n1944, 
            n1943, n1942, ram_s_131_6, n1941, ram_s_131_5, n1940, 
            ram_s_131_4, n1939, ram_s_131_3, n1938, ram_s_131_2, n1937, 
            ram_s_131_1, n1936, n1935, n1934, ram_s_130_6, n1933, 
            ram_s_130_5, n1932, ram_s_130_4, n1931, ram_s_130_3, n1930, 
            ram_s_130_2, n1929, ram_s_130_1, n1928, n1927, n1926, 
            ram_s_129_6, n1925, ram_s_129_5, n1924, ram_s_129_4, n1923, 
            ram_s_129_3, n1922, ram_s_129_2, n1921, ram_s_129_1, n1920, 
            n1919, n1918, ram_s_128_6, n1917, ram_s_128_5, n1916, 
            ram_s_128_4, n1915, ram_s_128_3, n1914, ram_s_128_2, n1913, 
            ram_s_128_1, n1912, n1543, ram_s_81_7, n1542, ram_s_81_6, 
            n1541, n1540, ram_s_81_4, n1539, ram_s_81_3, n1538, 
            ram_s_81_2, n1537, ram_s_81_1, n1536, ram_s_81_0, n1495, 
            n1494, ram_s_75_6, n1493, ram_s_75_5, n1492, n1491, 
            ram_s_75_3, n1490, n1489, ram_s_75_1, n1488, ram_s_75_0, 
            n1487, n1486, ram_s_74_6, n1485, ram_s_74_5, n1484, 
            n1483, ram_s_74_3, n1482, n1481, ram_s_74_1, n1480, 
            ram_s_74_0, n1479, n1478, ram_s_73_6, n1477, ram_s_73_5, 
            n1476, n1475, ram_s_73_3, n1474, n1473, ram_s_73_1, 
            n1472, ram_s_73_0, n1471, n1470, ram_s_72_6, n1469, 
            ram_s_72_5, n1468, n1467, ram_s_72_3, n1466, n1465, 
            ram_s_72_1, n1464, ram_s_72_0, n1463, ram_s_71_7, n1462, 
            ram_s_71_6, n1461, ram_s_71_5, n1460, n1459, n1458, 
            ram_s_71_2, n1457, ram_s_71_1, n1456, ram_s_71_0, n1455, 
            ram_s_70_7, n1454, ram_s_70_6, n1453, ram_s_70_5, n1452, 
            n1451, n1450, ram_s_70_2, n1449, ram_s_70_1, n1448, 
            ram_s_70_0, n1447, ram_s_69_7, n1446, ram_s_69_6, n1445, 
            ram_s_69_5, n1444, n1443, n1442, ram_s_69_2, n1441, 
            ram_s_69_1, n1440, ram_s_69_0, n1439, ram_s_68_7, n1438, 
            ram_s_68_6, n1437, ram_s_68_5, n1436, n1435, n1434, 
            ram_s_68_2, n1433, ram_s_68_1, n1432, ram_s_68_0, n1431, 
            ram_s_67_7, n1430, ram_s_67_6, n1429, ram_s_67_5, n1428, 
            n1427, ram_s_67_3, n1426, ram_s_67_2, n1425, ram_s_67_1, 
            n1424, n1423, ram_s_66_7, n1422, ram_s_66_6, n1421, 
            ram_s_66_5, n1420, n1419, ram_s_66_3, n1418, ram_s_66_2, 
            n1417, ram_s_66_1, n1416, n1415, ram_s_65_7, n1414, 
            ram_s_65_6, n1413, ram_s_65_5, n1412, n1411, ram_s_65_3, 
            n1410, ram_s_65_2, n1409, ram_s_65_1, n1408, n1407, 
            ram_s_64_7, n1406, ram_s_64_6, n1405, ram_s_64_5, n1404, 
            n1403, ram_s_64_3, n1402, ram_s_64_2, n1401, ram_s_64_1, 
            n1400, n1399, ram_s_63_7, n1398, ram_s_63_6, n1397, 
            ram_s_63_5, n1396, n1395, ram_s_63_3, n1394, ram_s_63_2, 
            n1393, ram_s_63_1, n1392, n1391, ram_s_62_7, n1390, 
            ram_s_62_6, n1389, ram_s_62_5, n1388, n1387, ram_s_62_3, 
            n1386, ram_s_62_2, n1385, ram_s_62_1, n1384, n1359, 
            ram_s_58_7, n1358, ram_s_58_6, n1357, n1356, ram_s_58_4, 
            n1355, ram_s_58_3, n1354, ram_s_58_2, n1353, ram_s_58_1, 
            n1352, n1351, ram_s_57_7, n1350, ram_s_57_6, n1349, 
            n1348, ram_s_57_4, n1347, ram_s_57_3, n1346, ram_s_57_2, 
            n1345, ram_s_57_1, n1344, n1271, ram_s_47_7, n1270, 
            ram_s_47_6, n1269, ram_s_47_5, n1268, ram_s_47_4, n1267, 
            ram_s_47_3, n1266, n1265, ram_s_47_1, n1264, ram_s_47_0, 
            n1255, ram_s_45_7, n1254, ram_s_45_6, n1253, ram_s_45_5, 
            n1252, ram_s_45_4, n1251, ram_s_45_3, n1250, n1249, 
            ram_s_45_1, n1248, ram_s_45_0, n1247, ram_s_44_7, n1246, 
            ram_s_44_6, n1245, ram_s_44_5, n1244, ram_s_44_4, n1243, 
            ram_s_44_3, n1242, n1241, ram_s_44_1, n1240, ram_s_44_0, 
            n1239, n1238, ram_s_43_6, n1237, ram_s_43_5, n1236, 
            ram_s_43_4, n1235, ram_s_43_3, n1234, n1233, n1232, 
            ram_s_43_0, n1215, n1214, ram_s_40_6, n1213, ram_s_40_5, 
            n1212, ram_s_40_4, n1211, ram_s_40_3, n1210, n1209, 
            n1208, ram_s_40_0, n1207, n1206, ram_s_39_6, n1205, 
            ram_s_39_5, n1204, ram_s_39_4, n1203, ram_s_39_3, n1202, 
            ram_s_39_2, n1201, ram_s_39_1, n1200, n1199, n1198, 
            ram_s_38_6, n1197, ram_s_38_5, n1196, ram_s_38_4, n1195, 
            ram_s_38_3, n1194, ram_s_38_2, n1193, ram_s_38_1, n1192, 
            n1191, n1190, ram_s_37_6, n1189, ram_s_37_5, n1188, 
            ram_s_37_4, n1187, ram_s_37_3, n1186, ram_s_37_2, n1185, 
            ram_s_37_1, n1184, n1183, n1182, ram_s_36_6, n1181, 
            ram_s_36_5, n1180, ram_s_36_4, n1179, ram_s_36_3, n1178, 
            ram_s_36_2, n1177, ram_s_36_1, n1176, n1175, n1174, 
            ram_s_35_6, n1173, ram_s_35_5, n1172, ram_s_35_4, n1171, 
            ram_s_35_3, n1170, n1169, n1168, ram_s_35_0, n1167, 
            n1166, ram_s_34_6, n1165, ram_s_34_5, n1164, ram_s_34_4, 
            n1163, ram_s_34_3, n1162, n1161, n1160, ram_s_34_0, 
            n1159, n1158, ram_s_33_6, n1157, ram_s_33_5, n1156, 
            ram_s_33_4, n1155, ram_s_33_3, n1154, n1153, n1152, 
            ram_s_33_0, n1151, n1150, ram_s_32_6, n1149, ram_s_32_5, 
            n1148, ram_s_32_4, n1147, ram_s_32_3, n1146, n1145, 
            n1144, ram_s_32_0, n1051, n1047, n1046, n1045, ram_s_0_2, 
            n1044, ram_s_12_3, n1043, n1042, ram_s_11_1, n1041, 
            n1040, ram_s_12_1, n1038, ram_s_11_4, n182, n1037, ram_s_12_4, 
            n54, n1036, ram_s_11_7, n183, n1035, n55, n1034, ram_s_12_7, 
            n184, n1033, ram_s_12_2, n56, n1032, ram_s_11_5, n185, 
            n1031, n57, n1030, ram_s_12_0, n186, n1029, ram_s_11_3, 
            n58, n187, n59, n188, n60, n189, n61, n190, n62, 
            n191, n63, n192, n1017, ram_s_0_3, n64, n1016, ram_s_0_4, 
            n193, n1015, ram_s_0_5, n65, n1014, ram_s_0_6, n194, 
            n1013, n66, n1012, n195, n1011, n67, n1010, ram_s_1_2, 
            n1009, ram_s_1_3, n1008, ram_s_1_4, n1007, ram_s_1_5, 
            n1006, ram_s_4_4, n1005, n1004, n1003, ram_s_5_0, n1002, 
            ram_s_4_6, n1001, ram_s_5_1, n998, ram_s_8_5, n997, 
            n996, n995, ram_s_7_4, n994, ram_s_7_1, n993, ram_s_6_6, 
            n992, ram_s_6_3, n989, n988, ram_s_8_3, n987, ram_s_8_0, 
            n986, n199, n985, ram_s_7_2, n71, n984, n200, n983, 
            ram_s_6_4, n72, n980, ram_s_8_7, n979, ram_s_8_4, n978, 
            ram_s_8_1, n977, ram_s_7_6, n976, ram_s_7_3, n975, ram_s_7_0, 
            n974, n973, ram_s_1_6, n972, n971, n970, n969, ram_s_2_2, 
            n968, ram_s_2_3, n967, ram_s_2_4, n966, ram_s_2_5, n965, 
            ram_s_2_6, n964, n963, n962, n961, ram_s_3_2, n960, 
            ram_s_3_3, n959, ram_s_3_4, n958, ram_s_3_5, n957, ram_s_14_7, 
            n952, ram_s_3_6, n950, n946, ram_s_4_0, n944, ram_s_4_1, 
            n941, ram_s_4_2, n940, ram_s_5_2, n939, ram_s_5_3, n935, 
            n934, ram_s_6_0, n933, ram_s_6_1, n932, ram_s_6_2, n931, 
            ram_s_5_6, n930, n927, ram_s_4_3, n926, n925, ram_s_13_3, 
            n924, ram_s_13_4, n923, n210, n82, n212, n84, n213, 
            n85, n214, n86, n217, n89, n218, n90, n219, n91, 
            n220, n92, n221, n93, n222, n94, n223, n95, n224, 
            n96, n225, n97, n918, ram_s_13_7, n917, ram_s_14_0, 
            n916, ram_s_14_1, spm_enable, n244, n116, n115, n243, 
            n245, n117, n246, n118, n48, n176, n249, n121, n250, 
            n122, n251, n123, n252, n124, n253, n125, n254, 
            n126, n255, n127, n256, n128, n257, n129, ram_s_14_2, 
            ram_s_13_2, ram_s_11_0, n911, n909, n908, ram_s_14_3, 
            n907, ram_s_13_1, n906, n904, ram_s_13_0, n901, ram_s_5_4, 
            n899);
    input [7:0]port_id;
    output ram_s_70_3;
    output ram_s_71_3;
    output ram_s_69_3;
    output ram_s_68_3;
    input \sx[7] ;
    input \sx[6] ;
    input \sx[5] ;
    input \sx[4] ;
    input \register_vector[10] ;
    output ram_s_34_7;
    output ram_s_35_7;
    output ram_s_33_7;
    output ram_s_32_7;
    input \register_vector[9] ;
    output ram_s_11_6;
    output ram_s_8_6;
    input \register_vector[11] ;
    output ram_s_62_4;
    output ram_s_63_4;
    output ram_s_2_7;
    output ram_s_3_7;
    output ram_s_1_7;
    output ram_s_0_7;
    output ram_s_66_4;
    output ram_s_67_4;
    output ram_s_65_4;
    output ram_s_64_4;
    input \register_vector[8] ;
    output ram_s_142_3;
    output ram_s_141_3;
    output ram_s_140_3;
    input CLK_3P3_MHZ_c;
    output ram_s_209_3;
    output ram_s_130_0;
    output ram_s_131_0;
    output ram_s_129_0;
    output ram_s_128_0;
    output ram_s_70_4;
    output ram_s_71_4;
    output ram_s_69_4;
    output ram_s_68_4;
    output ram_s_171_5;
    output ram_s_168_5;
    output ram_s_14_6;
    output ram_s_13_6;
    output ram_s_12_6;
    output ram_s_202_1;
    output ram_s_203_1;
    output ram_s_6_5;
    output ram_s_7_5;
    output ram_s_14_5;
    output ram_s_5_5;
    output ram_s_4_5;
    output ram_s_13_5;
    output ram_s_12_5;
    output ram_s_43_2;
    output ram_s_2_0;
    output ram_s_3_0;
    output ram_s_2_1;
    output ram_s_3_1;
    output ram_s_1_0;
    output ram_s_0_0;
    output ram_s_66_0;
    output ram_s_67_0;
    output ram_s_34_1;
    output ram_s_35_1;
    output ram_s_33_1;
    output ram_s_32_1;
    output ram_s_201_1;
    output ram_s_200_1;
    output ram_s_1_1;
    output ram_s_0_1;
    output ram_s_65_0;
    output ram_s_64_0;
    output ram_s_11_2;
    output ram_s_8_2;
    output ram_s_38_0;
    output ram_s_39_0;
    output ram_s_40_2;
    output ram_s_74_7;
    output ram_s_75_7;
    output ram_s_73_7;
    output ram_s_72_7;
    output ram_s_130_7;
    output ram_s_131_7;
    output ram_s_129_7;
    output ram_s_128_7;
    output ram_s_37_0;
    output ram_s_36_0;
    output ram_s_142_5;
    output ram_s_141_5;
    output ram_s_140_5;
    output ram_s_62_0;
    output ram_s_63_0;
    output ram_s_194_1;
    output ram_s_195_1;
    output ram_s_193_1;
    output ram_s_192_1;
    output ram_s_74_4;
    output ram_s_75_4;
    output ram_s_73_4;
    output ram_s_72_4;
    output ram_s_43_7;
    output ram_s_40_7;
    output ram_s_74_2;
    output ram_s_75_2;
    output ram_s_73_2;
    output ram_s_72_2;
    output ram_s_186_3;
    output ram_s_185_3;
    output ram_s_190_2;
    output ram_s_191_2;
    output ram_s_43_1;
    input [0:0]wea;
    output ram_s_40_1;
    output ram_s_6_7;
    output ram_s_7_7;
    output ram_s_134_0;
    output ram_s_135_0;
    output ram_s_5_7;
    output ram_s_4_7;
    output ram_s_133_0;
    output ram_s_132_0;
    output ram_s_34_2;
    output ram_s_35_2;
    output ram_s_58_5;
    output ram_s_58_0;
    output ram_s_57_0;
    output ram_s_139_0;
    output ram_s_136_0;
    output ram_s_190_5;
    output ram_s_191_5;
    output ram_s_57_5;
    output ram_s_33_2;
    output ram_s_32_2;
    output ram_s_142_7;
    output ram_s_141_7;
    output ram_s_140_7;
    output ram_s_81_5;
    output ram_s_190_1;
    output ram_s_191_1;
    output ram_s_139_1;
    output ram_s_136_1;
    output ram_s_38_7;
    output ram_s_39_7;
    output ram_s_37_7;
    output ram_s_36_7;
    input n893;
    output ram_s_14_4;
    output ram_s_190_7;
    output ram_s_191_7;
    output ram_s_47_2;
    output [7:0]spm_ram_data;
    output ram_s_45_2;
    output ram_s_44_2;
    output ram_s_134_5;
    output ram_s_135_5;
    output ram_s_133_5;
    output ram_s_132_5;
    input n2567;
    output ram_s_209_7;
    input n2566;
    output ram_s_209_6;
    input n2565;
    output ram_s_209_5;
    input n2564;
    output ram_s_209_4;
    input n2563;
    input n2562;
    output ram_s_209_2;
    input n2561;
    output ram_s_209_1;
    input n2560;
    output ram_s_209_0;
    input n2519;
    output ram_s_203_7;
    input n2518;
    output ram_s_203_6;
    input n2517;
    output ram_s_203_5;
    input n2516;
    output ram_s_203_4;
    input n2515;
    output ram_s_203_3;
    input n2514;
    output ram_s_203_2;
    input n2513;
    input n2512;
    output ram_s_203_0;
    input n2511;
    output ram_s_202_7;
    input n2510;
    output ram_s_202_6;
    input n2509;
    output ram_s_202_5;
    input n2508;
    output ram_s_202_4;
    input n2507;
    output ram_s_202_3;
    input n2506;
    output ram_s_202_2;
    input n2505;
    input n2504;
    output ram_s_202_0;
    input n2503;
    output ram_s_201_7;
    input n2502;
    output ram_s_201_6;
    input n2501;
    output ram_s_201_5;
    input n2500;
    output ram_s_201_4;
    input n2499;
    output ram_s_201_3;
    input n2498;
    output ram_s_201_2;
    input n2497;
    input n2496;
    output ram_s_201_0;
    input n2495;
    output ram_s_200_7;
    input n2494;
    output ram_s_200_6;
    input n2493;
    output ram_s_200_5;
    input n2492;
    output ram_s_200_4;
    input n2491;
    output ram_s_200_3;
    input n2490;
    output ram_s_200_2;
    input n2489;
    input n2488;
    output ram_s_200_0;
    input n2487;
    output ram_s_199_7;
    input n2486;
    output ram_s_199_6;
    input n2485;
    output ram_s_199_5;
    input n2484;
    output ram_s_199_4;
    input n2483;
    output ram_s_199_3;
    input n2482;
    output ram_s_199_2;
    input n2481;
    output ram_s_199_1;
    input n2480;
    output ram_s_199_0;
    input n2479;
    output ram_s_198_7;
    input n2478;
    output ram_s_198_6;
    input n2477;
    output ram_s_198_5;
    input n2476;
    output ram_s_198_4;
    input n2475;
    output ram_s_198_3;
    input n2474;
    output ram_s_198_2;
    input n2473;
    output ram_s_198_1;
    input n2472;
    output ram_s_198_0;
    input n2471;
    output ram_s_197_7;
    input n2470;
    output ram_s_197_6;
    input n2469;
    output ram_s_197_5;
    input n2468;
    output ram_s_197_4;
    input n2467;
    output ram_s_197_3;
    input n2466;
    output ram_s_197_2;
    input n2465;
    output ram_s_197_1;
    input n2464;
    output ram_s_197_0;
    input n2463;
    output ram_s_196_7;
    input n2462;
    output ram_s_196_6;
    input n2461;
    output ram_s_196_5;
    input n2460;
    output ram_s_196_4;
    input n2459;
    output ram_s_196_3;
    input n2458;
    output ram_s_196_2;
    input n2457;
    output ram_s_196_1;
    input n2456;
    output ram_s_196_0;
    input n2455;
    output ram_s_195_7;
    input n2454;
    output ram_s_195_6;
    input n2453;
    output ram_s_195_5;
    input n2452;
    output ram_s_195_4;
    input n2451;
    output ram_s_195_3;
    input n2450;
    output ram_s_195_2;
    input n2449;
    input n2448;
    output ram_s_195_0;
    input n2447;
    output ram_s_194_7;
    input n2446;
    output ram_s_194_6;
    input n2445;
    output ram_s_194_5;
    input n2444;
    output ram_s_194_4;
    input n2443;
    output ram_s_194_3;
    input n2442;
    output ram_s_194_2;
    input n2441;
    input n2440;
    output ram_s_194_0;
    input n2439;
    output ram_s_193_7;
    input n2438;
    output ram_s_193_6;
    input n2437;
    output ram_s_193_5;
    input n2436;
    output ram_s_193_4;
    input n2435;
    output ram_s_193_3;
    input n2434;
    output ram_s_193_2;
    input n2433;
    input n2432;
    output ram_s_193_0;
    input n2431;
    output ram_s_192_7;
    input n2430;
    output ram_s_192_6;
    input n2429;
    output ram_s_192_5;
    input n2428;
    output ram_s_192_4;
    input n2427;
    output ram_s_192_3;
    input n2426;
    output ram_s_192_2;
    input n2425;
    input n2424;
    output ram_s_192_0;
    input n2423;
    input n2422;
    output ram_s_191_6;
    input n2421;
    input n2420;
    output ram_s_191_4;
    input n2419;
    output ram_s_191_3;
    input n2418;
    input n2417;
    input n2416;
    output ram_s_191_0;
    input n2415;
    input n2414;
    output ram_s_190_6;
    input n2413;
    input n2412;
    output ram_s_190_4;
    input n2411;
    output ram_s_190_3;
    input n2410;
    input n2409;
    input n2408;
    output ram_s_190_0;
    input n2383;
    output ram_s_186_7;
    input n2382;
    output ram_s_186_6;
    input n2381;
    output ram_s_186_5;
    input n2380;
    output ram_s_186_4;
    input n2379;
    input n2378;
    output ram_s_186_2;
    input n2377;
    output ram_s_186_1;
    input n2376;
    output ram_s_186_0;
    input n2375;
    output ram_s_185_7;
    input n2374;
    output ram_s_185_6;
    input n2373;
    output ram_s_185_5;
    input n2372;
    output ram_s_185_4;
    input n2371;
    input n2370;
    output ram_s_185_2;
    input n2369;
    output ram_s_185_1;
    input n2368;
    output ram_s_185_0;
    input n2295;
    output ram_s_175_7;
    input n2294;
    output ram_s_175_6;
    input n2293;
    output ram_s_175_5;
    input n2292;
    output ram_s_175_4;
    input n2291;
    output ram_s_175_3;
    input n2290;
    output ram_s_175_2;
    input n2289;
    output ram_s_175_1;
    input n2288;
    output ram_s_175_0;
    input n2279;
    output ram_s_173_7;
    input n2278;
    output ram_s_173_6;
    input n2277;
    output ram_s_173_5;
    input n2276;
    output ram_s_173_4;
    input n2275;
    output ram_s_173_3;
    input n2274;
    output ram_s_173_2;
    input n2273;
    output ram_s_173_1;
    input n2272;
    output ram_s_173_0;
    input n2271;
    output ram_s_172_7;
    input n2270;
    output ram_s_172_6;
    input n2269;
    output ram_s_172_5;
    input n2268;
    output ram_s_172_4;
    input n2267;
    output ram_s_172_3;
    input n2266;
    output ram_s_172_2;
    input n2265;
    output ram_s_172_1;
    input n2264;
    output ram_s_172_0;
    input n2263;
    output ram_s_171_7;
    input n2262;
    output ram_s_171_6;
    input n2261;
    input n2260;
    output ram_s_171_4;
    input n2259;
    output ram_s_171_3;
    input n2258;
    output ram_s_171_2;
    input n2257;
    output ram_s_171_1;
    input n2256;
    output ram_s_171_0;
    input n2239;
    output ram_s_168_7;
    input n2238;
    output ram_s_168_6;
    input n2237;
    input n2236;
    output ram_s_168_4;
    input n2235;
    output ram_s_168_3;
    input n2234;
    output ram_s_168_2;
    input n2233;
    output ram_s_168_1;
    input n2232;
    output ram_s_168_0;
    input n2231;
    output ram_s_167_7;
    input n2230;
    output ram_s_167_6;
    input n2229;
    output ram_s_167_5;
    input n2228;
    output ram_s_167_4;
    input n2227;
    output ram_s_167_3;
    input n2226;
    output ram_s_167_2;
    input n2225;
    output ram_s_167_1;
    input n2224;
    output ram_s_167_0;
    input n2223;
    output ram_s_166_7;
    input n2222;
    output ram_s_166_6;
    input n2221;
    output ram_s_166_5;
    input n2220;
    output ram_s_166_4;
    input n2219;
    output ram_s_166_3;
    input n2218;
    output ram_s_166_2;
    input n2217;
    output ram_s_166_1;
    input n2216;
    output ram_s_166_0;
    input n2215;
    output ram_s_165_7;
    input n2214;
    output ram_s_165_6;
    input n2213;
    output ram_s_165_5;
    input n2212;
    output ram_s_165_4;
    input n2211;
    output ram_s_165_3;
    input n2210;
    output ram_s_165_2;
    input n2209;
    output ram_s_165_1;
    input n2208;
    output ram_s_165_0;
    input n2207;
    output ram_s_164_7;
    input n2206;
    output ram_s_164_6;
    input n2205;
    output ram_s_164_5;
    input n2204;
    output ram_s_164_4;
    input n2203;
    output ram_s_164_3;
    input n2202;
    output ram_s_164_2;
    input n2201;
    output ram_s_164_1;
    input n2200;
    output ram_s_164_0;
    input n2199;
    output ram_s_163_7;
    input n2198;
    output ram_s_163_6;
    input n2197;
    output ram_s_163_5;
    input n2196;
    output ram_s_163_4;
    input n2195;
    output ram_s_163_3;
    input n2194;
    output ram_s_163_2;
    input n2193;
    output ram_s_163_1;
    input n2192;
    output ram_s_163_0;
    input n2191;
    output ram_s_162_7;
    input n2190;
    output ram_s_162_6;
    input n2189;
    output ram_s_162_5;
    input n2188;
    output ram_s_162_4;
    input n2187;
    output ram_s_162_3;
    input n2186;
    output ram_s_162_2;
    input n2185;
    output ram_s_162_1;
    input n2184;
    output ram_s_162_0;
    input n2183;
    output ram_s_161_7;
    input n2182;
    output ram_s_161_6;
    input n2181;
    output ram_s_161_5;
    input n2180;
    output ram_s_161_4;
    input n2179;
    output ram_s_161_3;
    input n2178;
    output ram_s_161_2;
    input n2177;
    output ram_s_161_1;
    input n2176;
    output ram_s_161_0;
    input n2175;
    output ram_s_160_7;
    input n2174;
    output ram_s_160_6;
    input n2173;
    output ram_s_160_5;
    input n2172;
    output ram_s_160_4;
    input n2171;
    output ram_s_160_3;
    input n2170;
    output ram_s_160_2;
    input n2169;
    output ram_s_160_1;
    input n2168;
    output ram_s_160_0;
    input n2031;
    input n2030;
    output ram_s_142_6;
    input n2029;
    input n2028;
    output ram_s_142_4;
    input n2027;
    input n2026;
    output ram_s_142_2;
    input n2025;
    output ram_s_142_1;
    input n2024;
    output ram_s_142_0;
    input n2023;
    input n2022;
    output ram_s_141_6;
    input n2021;
    input n2020;
    output ram_s_141_4;
    input n2019;
    input n2018;
    output ram_s_141_2;
    input n2017;
    output ram_s_141_1;
    input n2016;
    output ram_s_141_0;
    input n2015;
    input n2014;
    output ram_s_140_6;
    input n2013;
    input n2012;
    output ram_s_140_4;
    input n2011;
    input n2010;
    output ram_s_140_2;
    input n2009;
    output ram_s_140_1;
    input n2008;
    output ram_s_140_0;
    input n2007;
    output ram_s_139_7;
    input n2006;
    output ram_s_139_6;
    input n2005;
    output ram_s_139_5;
    input n2004;
    output ram_s_139_4;
    input n2003;
    output ram_s_139_3;
    input n2002;
    output ram_s_139_2;
    input n2001;
    input n2000;
    input n1983;
    output ram_s_136_7;
    input n1982;
    output ram_s_136_6;
    input n1981;
    output ram_s_136_5;
    input n1980;
    output ram_s_136_4;
    input n1979;
    output ram_s_136_3;
    input n1978;
    output ram_s_136_2;
    input n1977;
    input n1976;
    input n1975;
    output ram_s_135_7;
    input n1974;
    output ram_s_135_6;
    input n1973;
    input n1972;
    output ram_s_135_4;
    input n1971;
    output ram_s_135_3;
    input n1970;
    output ram_s_135_2;
    input n1969;
    output ram_s_135_1;
    input n1968;
    input n1967;
    output ram_s_134_7;
    input n1966;
    output ram_s_134_6;
    input n1965;
    input n1964;
    output ram_s_134_4;
    input n1963;
    output ram_s_134_3;
    input n1962;
    output ram_s_134_2;
    input n1961;
    output ram_s_134_1;
    input n1960;
    input n1959;
    output ram_s_133_7;
    input n1958;
    output ram_s_133_6;
    input n1957;
    input n1956;
    output ram_s_133_4;
    input n1955;
    output ram_s_133_3;
    input n1954;
    output ram_s_133_2;
    input n1953;
    output ram_s_133_1;
    input n1952;
    input n1951;
    output ram_s_132_7;
    input n1950;
    output ram_s_132_6;
    input n1949;
    input n1948;
    output ram_s_132_4;
    input n1947;
    output ram_s_132_3;
    input n1946;
    output ram_s_132_2;
    input n1945;
    output ram_s_132_1;
    input n1944;
    input n1943;
    input n1942;
    output ram_s_131_6;
    input n1941;
    output ram_s_131_5;
    input n1940;
    output ram_s_131_4;
    input n1939;
    output ram_s_131_3;
    input n1938;
    output ram_s_131_2;
    input n1937;
    output ram_s_131_1;
    input n1936;
    input n1935;
    input n1934;
    output ram_s_130_6;
    input n1933;
    output ram_s_130_5;
    input n1932;
    output ram_s_130_4;
    input n1931;
    output ram_s_130_3;
    input n1930;
    output ram_s_130_2;
    input n1929;
    output ram_s_130_1;
    input n1928;
    input n1927;
    input n1926;
    output ram_s_129_6;
    input n1925;
    output ram_s_129_5;
    input n1924;
    output ram_s_129_4;
    input n1923;
    output ram_s_129_3;
    input n1922;
    output ram_s_129_2;
    input n1921;
    output ram_s_129_1;
    input n1920;
    input n1919;
    input n1918;
    output ram_s_128_6;
    input n1917;
    output ram_s_128_5;
    input n1916;
    output ram_s_128_4;
    input n1915;
    output ram_s_128_3;
    input n1914;
    output ram_s_128_2;
    input n1913;
    output ram_s_128_1;
    input n1912;
    input n1543;
    output ram_s_81_7;
    input n1542;
    output ram_s_81_6;
    input n1541;
    input n1540;
    output ram_s_81_4;
    input n1539;
    output ram_s_81_3;
    input n1538;
    output ram_s_81_2;
    input n1537;
    output ram_s_81_1;
    input n1536;
    output ram_s_81_0;
    input n1495;
    input n1494;
    output ram_s_75_6;
    input n1493;
    output ram_s_75_5;
    input n1492;
    input n1491;
    output ram_s_75_3;
    input n1490;
    input n1489;
    output ram_s_75_1;
    input n1488;
    output ram_s_75_0;
    input n1487;
    input n1486;
    output ram_s_74_6;
    input n1485;
    output ram_s_74_5;
    input n1484;
    input n1483;
    output ram_s_74_3;
    input n1482;
    input n1481;
    output ram_s_74_1;
    input n1480;
    output ram_s_74_0;
    input n1479;
    input n1478;
    output ram_s_73_6;
    input n1477;
    output ram_s_73_5;
    input n1476;
    input n1475;
    output ram_s_73_3;
    input n1474;
    input n1473;
    output ram_s_73_1;
    input n1472;
    output ram_s_73_0;
    input n1471;
    input n1470;
    output ram_s_72_6;
    input n1469;
    output ram_s_72_5;
    input n1468;
    input n1467;
    output ram_s_72_3;
    input n1466;
    input n1465;
    output ram_s_72_1;
    input n1464;
    output ram_s_72_0;
    input n1463;
    output ram_s_71_7;
    input n1462;
    output ram_s_71_6;
    input n1461;
    output ram_s_71_5;
    input n1460;
    input n1459;
    input n1458;
    output ram_s_71_2;
    input n1457;
    output ram_s_71_1;
    input n1456;
    output ram_s_71_0;
    input n1455;
    output ram_s_70_7;
    input n1454;
    output ram_s_70_6;
    input n1453;
    output ram_s_70_5;
    input n1452;
    input n1451;
    input n1450;
    output ram_s_70_2;
    input n1449;
    output ram_s_70_1;
    input n1448;
    output ram_s_70_0;
    input n1447;
    output ram_s_69_7;
    input n1446;
    output ram_s_69_6;
    input n1445;
    output ram_s_69_5;
    input n1444;
    input n1443;
    input n1442;
    output ram_s_69_2;
    input n1441;
    output ram_s_69_1;
    input n1440;
    output ram_s_69_0;
    input n1439;
    output ram_s_68_7;
    input n1438;
    output ram_s_68_6;
    input n1437;
    output ram_s_68_5;
    input n1436;
    input n1435;
    input n1434;
    output ram_s_68_2;
    input n1433;
    output ram_s_68_1;
    input n1432;
    output ram_s_68_0;
    input n1431;
    output ram_s_67_7;
    input n1430;
    output ram_s_67_6;
    input n1429;
    output ram_s_67_5;
    input n1428;
    input n1427;
    output ram_s_67_3;
    input n1426;
    output ram_s_67_2;
    input n1425;
    output ram_s_67_1;
    input n1424;
    input n1423;
    output ram_s_66_7;
    input n1422;
    output ram_s_66_6;
    input n1421;
    output ram_s_66_5;
    input n1420;
    input n1419;
    output ram_s_66_3;
    input n1418;
    output ram_s_66_2;
    input n1417;
    output ram_s_66_1;
    input n1416;
    input n1415;
    output ram_s_65_7;
    input n1414;
    output ram_s_65_6;
    input n1413;
    output ram_s_65_5;
    input n1412;
    input n1411;
    output ram_s_65_3;
    input n1410;
    output ram_s_65_2;
    input n1409;
    output ram_s_65_1;
    input n1408;
    input n1407;
    output ram_s_64_7;
    input n1406;
    output ram_s_64_6;
    input n1405;
    output ram_s_64_5;
    input n1404;
    input n1403;
    output ram_s_64_3;
    input n1402;
    output ram_s_64_2;
    input n1401;
    output ram_s_64_1;
    input n1400;
    input n1399;
    output ram_s_63_7;
    input n1398;
    output ram_s_63_6;
    input n1397;
    output ram_s_63_5;
    input n1396;
    input n1395;
    output ram_s_63_3;
    input n1394;
    output ram_s_63_2;
    input n1393;
    output ram_s_63_1;
    input n1392;
    input n1391;
    output ram_s_62_7;
    input n1390;
    output ram_s_62_6;
    input n1389;
    output ram_s_62_5;
    input n1388;
    input n1387;
    output ram_s_62_3;
    input n1386;
    output ram_s_62_2;
    input n1385;
    output ram_s_62_1;
    input n1384;
    input n1359;
    output ram_s_58_7;
    input n1358;
    output ram_s_58_6;
    input n1357;
    input n1356;
    output ram_s_58_4;
    input n1355;
    output ram_s_58_3;
    input n1354;
    output ram_s_58_2;
    input n1353;
    output ram_s_58_1;
    input n1352;
    input n1351;
    output ram_s_57_7;
    input n1350;
    output ram_s_57_6;
    input n1349;
    input n1348;
    output ram_s_57_4;
    input n1347;
    output ram_s_57_3;
    input n1346;
    output ram_s_57_2;
    input n1345;
    output ram_s_57_1;
    input n1344;
    input n1271;
    output ram_s_47_7;
    input n1270;
    output ram_s_47_6;
    input n1269;
    output ram_s_47_5;
    input n1268;
    output ram_s_47_4;
    input n1267;
    output ram_s_47_3;
    input n1266;
    input n1265;
    output ram_s_47_1;
    input n1264;
    output ram_s_47_0;
    input n1255;
    output ram_s_45_7;
    input n1254;
    output ram_s_45_6;
    input n1253;
    output ram_s_45_5;
    input n1252;
    output ram_s_45_4;
    input n1251;
    output ram_s_45_3;
    input n1250;
    input n1249;
    output ram_s_45_1;
    input n1248;
    output ram_s_45_0;
    input n1247;
    output ram_s_44_7;
    input n1246;
    output ram_s_44_6;
    input n1245;
    output ram_s_44_5;
    input n1244;
    output ram_s_44_4;
    input n1243;
    output ram_s_44_3;
    input n1242;
    input n1241;
    output ram_s_44_1;
    input n1240;
    output ram_s_44_0;
    input n1239;
    input n1238;
    output ram_s_43_6;
    input n1237;
    output ram_s_43_5;
    input n1236;
    output ram_s_43_4;
    input n1235;
    output ram_s_43_3;
    input n1234;
    input n1233;
    input n1232;
    output ram_s_43_0;
    input n1215;
    input n1214;
    output ram_s_40_6;
    input n1213;
    output ram_s_40_5;
    input n1212;
    output ram_s_40_4;
    input n1211;
    output ram_s_40_3;
    input n1210;
    input n1209;
    input n1208;
    output ram_s_40_0;
    input n1207;
    input n1206;
    output ram_s_39_6;
    input n1205;
    output ram_s_39_5;
    input n1204;
    output ram_s_39_4;
    input n1203;
    output ram_s_39_3;
    input n1202;
    output ram_s_39_2;
    input n1201;
    output ram_s_39_1;
    input n1200;
    input n1199;
    input n1198;
    output ram_s_38_6;
    input n1197;
    output ram_s_38_5;
    input n1196;
    output ram_s_38_4;
    input n1195;
    output ram_s_38_3;
    input n1194;
    output ram_s_38_2;
    input n1193;
    output ram_s_38_1;
    input n1192;
    input n1191;
    input n1190;
    output ram_s_37_6;
    input n1189;
    output ram_s_37_5;
    input n1188;
    output ram_s_37_4;
    input n1187;
    output ram_s_37_3;
    input n1186;
    output ram_s_37_2;
    input n1185;
    output ram_s_37_1;
    input n1184;
    input n1183;
    input n1182;
    output ram_s_36_6;
    input n1181;
    output ram_s_36_5;
    input n1180;
    output ram_s_36_4;
    input n1179;
    output ram_s_36_3;
    input n1178;
    output ram_s_36_2;
    input n1177;
    output ram_s_36_1;
    input n1176;
    input n1175;
    input n1174;
    output ram_s_35_6;
    input n1173;
    output ram_s_35_5;
    input n1172;
    output ram_s_35_4;
    input n1171;
    output ram_s_35_3;
    input n1170;
    input n1169;
    input n1168;
    output ram_s_35_0;
    input n1167;
    input n1166;
    output ram_s_34_6;
    input n1165;
    output ram_s_34_5;
    input n1164;
    output ram_s_34_4;
    input n1163;
    output ram_s_34_3;
    input n1162;
    input n1161;
    input n1160;
    output ram_s_34_0;
    input n1159;
    input n1158;
    output ram_s_33_6;
    input n1157;
    output ram_s_33_5;
    input n1156;
    output ram_s_33_4;
    input n1155;
    output ram_s_33_3;
    input n1154;
    input n1153;
    input n1152;
    output ram_s_33_0;
    input n1151;
    input n1150;
    output ram_s_32_6;
    input n1149;
    output ram_s_32_5;
    input n1148;
    output ram_s_32_4;
    input n1147;
    output ram_s_32_3;
    input n1146;
    input n1145;
    input n1144;
    output ram_s_32_0;
    input n1051;
    input n1047;
    input n1046;
    input n1045;
    output ram_s_0_2;
    input n1044;
    output ram_s_12_3;
    input n1043;
    input n1042;
    output ram_s_11_1;
    input n1041;
    input n1040;
    output ram_s_12_1;
    input n1038;
    output ram_s_11_4;
    output n182;
    input n1037;
    output ram_s_12_4;
    output n54;
    input n1036;
    output ram_s_11_7;
    output n183;
    input n1035;
    output n55;
    input n1034;
    output ram_s_12_7;
    output n184;
    input n1033;
    output ram_s_12_2;
    output n56;
    input n1032;
    output ram_s_11_5;
    output n185;
    input n1031;
    output n57;
    input n1030;
    output ram_s_12_0;
    output n186;
    input n1029;
    output ram_s_11_3;
    output n58;
    output n187;
    output n59;
    output n188;
    output n60;
    output n189;
    output n61;
    output n190;
    output n62;
    output n191;
    output n63;
    output n192;
    input n1017;
    output ram_s_0_3;
    output n64;
    input n1016;
    output ram_s_0_4;
    output n193;
    input n1015;
    output ram_s_0_5;
    output n65;
    input n1014;
    output ram_s_0_6;
    output n194;
    input n1013;
    output n66;
    input n1012;
    output n195;
    input n1011;
    output n67;
    input n1010;
    output ram_s_1_2;
    input n1009;
    output ram_s_1_3;
    input n1008;
    output ram_s_1_4;
    input n1007;
    output ram_s_1_5;
    input n1006;
    output ram_s_4_4;
    input n1005;
    input n1004;
    input n1003;
    output ram_s_5_0;
    input n1002;
    output ram_s_4_6;
    input n1001;
    output ram_s_5_1;
    input n998;
    output ram_s_8_5;
    input n997;
    input n996;
    input n995;
    output ram_s_7_4;
    input n994;
    output ram_s_7_1;
    input n993;
    output ram_s_6_6;
    input n992;
    output ram_s_6_3;
    input n989;
    input n988;
    output ram_s_8_3;
    input n987;
    output ram_s_8_0;
    input n986;
    output n199;
    input n985;
    output ram_s_7_2;
    output n71;
    input n984;
    output n200;
    input n983;
    output ram_s_6_4;
    output n72;
    input n980;
    output ram_s_8_7;
    input n979;
    output ram_s_8_4;
    input n978;
    output ram_s_8_1;
    input n977;
    output ram_s_7_6;
    input n976;
    output ram_s_7_3;
    input n975;
    output ram_s_7_0;
    input n974;
    input n973;
    output ram_s_1_6;
    input n972;
    input n971;
    input n970;
    input n969;
    output ram_s_2_2;
    input n968;
    output ram_s_2_3;
    input n967;
    output ram_s_2_4;
    input n966;
    output ram_s_2_5;
    input n965;
    output ram_s_2_6;
    input n964;
    input n963;
    input n962;
    input n961;
    output ram_s_3_2;
    input n960;
    output ram_s_3_3;
    input n959;
    output ram_s_3_4;
    input n958;
    output ram_s_3_5;
    input n957;
    output ram_s_14_7;
    input n952;
    output ram_s_3_6;
    input n950;
    input n946;
    output ram_s_4_0;
    input n944;
    output ram_s_4_1;
    input n941;
    output ram_s_4_2;
    input n940;
    output ram_s_5_2;
    input n939;
    output ram_s_5_3;
    input n935;
    input n934;
    output ram_s_6_0;
    input n933;
    output ram_s_6_1;
    input n932;
    output ram_s_6_2;
    input n931;
    output ram_s_5_6;
    input n930;
    input n927;
    output ram_s_4_3;
    input n926;
    input n925;
    output ram_s_13_3;
    input n924;
    output ram_s_13_4;
    input n923;
    output n210;
    output n82;
    output n212;
    output n84;
    output n213;
    output n85;
    output n214;
    output n86;
    output n217;
    output n89;
    output n218;
    output n90;
    output n219;
    output n91;
    output n220;
    output n92;
    output n221;
    output n93;
    output n222;
    output n94;
    output n223;
    output n95;
    output n224;
    output n96;
    output n225;
    output n97;
    input n918;
    output ram_s_13_7;
    input n917;
    output ram_s_14_0;
    input n916;
    output ram_s_14_1;
    input spm_enable;
    output n244;
    output n116;
    output n115;
    output n243;
    output n245;
    output n117;
    output n246;
    output n118;
    output n48;
    output n176;
    output n249;
    output n121;
    output n250;
    output n122;
    output n251;
    output n123;
    output n252;
    output n124;
    output n253;
    output n125;
    output n254;
    output n126;
    output n255;
    output n127;
    output n256;
    output n128;
    output n257;
    output n129;
    output ram_s_14_2;
    output ram_s_13_2;
    output ram_s_11_0;
    input n911;
    input n909;
    input n908;
    output ram_s_14_3;
    input n907;
    output ram_s_13_1;
    input n906;
    input n904;
    output ram_s_13_0;
    input n901;
    output ram_s_5_4;
    input n899;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    wire n13199, n9038, ram_s_154_6, ram_s_155_6, n13193, ram_s_153_6, 
        ram_s_152_6, n13196, ram_s_254_0, ram_s_255_0, n13187, ram_s_253_0, 
        ram_s_252_0, n13190, n177, ram_s_85_7, n1575, n237, ram_s_115_7, 
        n1815, ram_s_85_6, n1574, ram_s_115_6, n1814, ram_s_115_5, 
        n1813, ram_s_115_4, n1812, n161, ram_s_77_2, n1506, n13181, 
        n13184, n159, ram_s_76_1, n1497, ram_s_10_6, n13175, ram_s_9_6, 
        n9044, ram_s_85_5, n1573, ram_s_115_3, n1811, n9495, n9496, 
        n13169, n9484, n9483, n13172, ram_s_250_2, ram_s_251_2, 
        n13163, ram_s_115_2, n1810, ram_s_249_2, ram_s_248_2, n13166, 
        ram_s_85_4, n1572, ram_s_126_0, ram_s_127_0, n13157, ram_s_115_1, 
        n1809, ram_s_125_0, ram_s_124_0, n9047, n13004, n9451, n13151, 
        n9445, n12992, n13154, n10025, n10043, n13145, n10004, 
        n9995, n13139, ram_s_61_4, ram_s_60_4, n9671, n13133, n13136, 
        n13127, n9674, n12260, n12194, n13121, n12272, n12356, 
        n13124, ram_s_115_0, n1808, ram_s_254_2, ram_s_255_2, n13115, 
        ram_s_253_2, ram_s_252_2, n13118, n225_c, ram_s_237_7, n2791, 
        n10604, n10610, n13109, n10589, n10586, n10805, ram_s_246_5, 
        ram_s_247_5, n13103, ram_s_245_5, ram_s_244_5, n10418, ram_s_143_3, 
        n13097, n9680, ram_s_237_6, n2790, ram_s_158_6, ram_s_159_6, 
        n13091, ram_s_157_6, ram_s_156_6, n13094, ram_s_237_5, n2789, 
        ram_s_237_4, n2788, ram_s_178_2, ram_s_179_2, n13085, ram_s_177_2, 
        ram_s_176_2, n13088, n9336, n9337, n13079, ram_s_237_3, 
        n2787, n9328, n9327, n13082, ram_s_237_2, n2786, n898, 
        ram_s_10_2, ram_s_85_3, n1571, ram_s_210_3, ram_s_211_3, n11225, 
        ram_s_237_1, n2785, ram_s_208_3, n11228, ram_s_237_0, n2784, 
        ram_s_85_2, n1570, n13073, ram_s_85_1, n1569, n235, ram_s_114_7, 
        n1807, ram_s_114_6, n1806, n9053, ram_s_114_5, n1805, ram_s_114_4, 
        n1804, n13067, ram_s_114_3, n1803, ram_s_30_1, ram_s_31_1, 
        n12137, n9686, ram_s_29_1, ram_s_28_1, n12140, ram_s_170_5, 
        n13061, ram_s_169_5, n9347, n9312, n9313, n13055, n9304, 
        n9303, n13058, ram_s_15_6, n13049, n9056, n9282, n9283, 
        n13043, n9262, n9261, n13046, ram_s_114_2, n1802, ram_s_114_1, 
        n1801, n11219, n12359, ram_s_15_5, n11939, n10469, n9966, 
        n9967, n11513, n11006, ram_s_114_0, n1800, n9955, n9954, 
        n11516, ram_s_42_2, n11747, n12353, n13031, n223_c, ram_s_236_7, 
        n2783, ram_s_236_6, n2782, ram_s_236_5, n2781, n11507, n12125, 
        n9764, n11606, n11933, n12128, n9758, n9740, n11009, n11222, 
        ram_s_236_4, n2780, n13034, ram_s_236_3, n2779, n11510, 
        n13025, ram_s_9_2, n10808, ram_s_146_7, ram_s_147_7, n11213, 
        n11501, ram_s_236_2, n2778, n10278, n10279, n12347, ram_s_178_6, 
        ram_s_179_6, n12119, ram_s_236_1, n2777, ram_s_41_2, n11750, 
        ram_s_177_6, ram_s_176_6, n12122, n13019, n10264, n10263, 
        n10882, ram_s_236_0, n2776, ram_s_113_2, ram_s_112_2, n13022, 
        ram_s_145_7, ram_s_144_7, n11216, n12032, n11978, n13013, 
        n11678, n9116, n12113, n12068, n12110, n13016, n11186, 
        n9809, n11921, n11486, n11600, n11015, n13007, n9017, 
        n12116, n13010, n12341, n9240, n9241, n13001, ram_s_77_1, 
        n1505, n12344, ram_s_18_0, ram_s_19_0, n12107, ram_s_85_0, 
        n1568, n173, ram_s_211_7, n2583, n233, ram_s_113_7, n1799, 
        n11504, ram_s_113_6, n1798, ram_s_113_5, n1797, ram_s_211_6, 
        n2582, ram_s_211_5, n2581, ram_s_113_4, n1796, ram_s_143_5, 
        n11735, ram_s_113_3, n1795, ram_s_17_0, ram_s_16_0, n11738, 
        n1794, ram_s_113_1, n1793, n9232, n9231, ram_s_30_5, ram_s_31_5, 
        n12335, ram_s_113_0, n1792, n221_c, ram_s_235_7, n2775, 
        n11729, ram_s_211_4, n2580, n11585, ram_s_235_6, n2774, 
        ram_s_29_5, ram_s_28_5, n9752, n2579, n11909, ram_s_61_0, 
        ram_s_60_0, n11732, ram_s_235_5, n2773, ram_s_211_2, n2578, 
        n11588, ram_s_235_4, n2772, ram_s_77_0, n1504, n9207, n9208, 
        n12989, n9196, n9195, n9023, n9008, n11912, n12983, n9692, 
        ram_s_42_7, n11723, ram_s_41_7, n11726, n9264, n9265, n12971, 
        ram_s_235_3, n2771, n11207, ram_s_235_2, n2770, n11210, 
        ram_s_235_1, n2769, ram_s_235_0, n2768, n9794, n9818, n11201, 
        ram_s_86_7, ram_s_87_7, n11579, n9746, n9725, n11204, n219_c, 
        ram_s_234_7, n2767, n165, ram_s_207_7, n2551, ram_s_234_6, 
        n2766, ram_s_234_5, n2765, n9253, n9252, n12974, ram_s_211_1, 
        n2577, ram_s_234_4, n2764, ram_s_187_3, n12965, ram_s_184_3, 
        n12968, n9171, n9172, n12959, n9163, n9162, n12962, ram_s_76_0, 
        n1496, ram_s_207_6, n2550, ram_s_206_7, n12095, ram_s_84_7, 
        n11582, n10634, n10649, n12953, n10625, n10622, n10811, 
        ram_s_214_7, ram_s_215_7, n11717, n12329, ram_s_205_7, ram_s_204_7, 
        n10499, ram_s_213_7, ram_s_212_7, n10532, ram_s_234_3, n2763, 
        ram_s_42_1, n11573, ram_s_234_2, n2762, ram_s_211_0, n2576, 
        n45, n174, ram_s_234_1, n2761, ram_s_234_0, n2760, n231, 
        ram_s_112_7, n1791, ram_s_112_6, n1790, ram_s_112_5, n1789, 
        ram_s_112_4, n1788, ram_s_41_1, n11576, ram_s_112_3, n1787, 
        n1786, ram_s_112_1, n1785, ram_s_112_0, n1784, n217_c, ram_s_233_7, 
        n2759, ram_s_233_6, n2758, ram_s_233_5, n2757, ram_s_233_4, 
        n2756, n11711, ram_s_233_3, n2755, n12947, n11714, n9065, 
        ram_s_189_2, ram_s_188_2, n12332, n12089, ram_s_233_2, n2754, 
        ram_s_233_1, n2753, n175, n1567, ram_s_84_6, n1566, ram_s_84_5, 
        n1565, ram_s_84_4, n1564, ram_s_84_3, n1563, ram_s_84_2, 
        n1562, ram_s_84_1, n1561, ram_s_84_0, n1560, n9855, n9856, 
        n12941, ram_s_233_0, n2752, n9814, n9813, n10813, n229, 
        ram_s_111_7, n1783, ram_s_59_5, n11705, n9141, n9142, n12935, 
        n171, ram_s_210_7, n2575, ram_s_111_6, n1782, n9127, n9126, 
        n12938, ram_s_182_2, ram_s_183_2, n12929, ram_s_181_2, ram_s_180_2, 
        n12932, ram_s_111_5, n1781, ram_s_111_4, n1780, ram_s_111_3, 
        n1779, ram_s_111_2, n1778, ram_s_111_1, n1777, ram_s_111_0, 
        n1776, ram_s_50_0, ram_s_51_0, n11195, n10541, n11252, n11567, 
        ram_s_59_0, n12917, ram_s_56_0, n8906, ram_s_94_5, ram_s_95_5, 
        n12911, ram_s_93_5, ram_s_92_5, n12914, n12698, n12905, 
        n10796, n10772, n12908, ram_s_138_0, n12899, ram_s_137_0, 
        n9068, n9135, n9136, n12893, ram_s_210_6, n2574, n215, 
        ram_s_232_7, n2751, ram_s_232_6, n2750, n10517, n11570, 
        n9061, n9060, n10816, n12887, ram_s_189_5, ram_s_188_5, 
        n9701, n11456, n11288, n12881, n11774, n12884, ram_s_250_4, 
        ram_s_251_4, n12875, ram_s_232_5, n2749, ram_s_232_4, n2748, 
        ram_s_249_4, ram_s_248_4, n12878, n12869, ram_s_56_5, n11708, 
        n12092, n9872, n9881, n11891, ram_s_143_7, n11561, ram_s_210_5, 
        n2573, n9863, n9854, n11033, n11966, n11198, n12872, n11564, 
        ram_s_110_3, n12323, ram_s_94_6, ram_s_95_6, n11699, ram_s_109_3, 
        ram_s_108_3, n9395, ram_s_93_6, ram_s_92_6, n11702, ram_s_82_5, 
        ram_s_83_5, n12863, ram_s_80_5, n12866, ram_s_232_3, n2747, 
        ram_s_158_1, ram_s_159_1, n12317, ram_s_157_1, ram_s_156_1, 
        n12320, n11693, ram_s_49_0, ram_s_48_0, n897, ram_s_138_1, 
        n12857, n9662, n11885, n9999, n10000, n11189, n9644, n9635, 
        n11888, ram_s_137_1, n12860, n896, ram_s_10_0, n895, ram_s_10_3, 
        n12851, n894, ram_s_10_1, n12854, n9991, n9990, n11192, 
        ram_s_232_2, n2746, ram_s_250_6, ram_s_251_6, n12845, n892, 
        ram_s_21_3, ram_s_249_6, ram_s_248_6, n12848, n891, n890, 
        ram_s_17_1, ram_s_232_1, n2745, ram_s_78_4, ram_s_79_4, n12839, 
        n889, ram_s_17_2, ram_s_232_0, n2744, ram_s_77_4, ram_s_76_4, 
        n9707, ram_s_210_4, n2572, n888, ram_s_17_3, n12833, ram_s_189_7, 
        ram_s_188_7, n10427, ram_s_118_4, ram_s_119_4, n11483, ram_s_122_4, 
        ram_s_123_4, n11183, ram_s_117_4, ram_s_116_4, ram_s_46_2, 
        n11477, n227, ram_s_110_7, n1775, n887, ram_s_17_4, n886, 
        ram_s_10_4, n885, ram_s_17_5, ram_s_110_6, n1774, n11480, 
        ram_s_110_5, n1773, ram_s_110_4, n1772, n1771, ram_s_110_2, 
        n1770, ram_s_110_1, n1769, ram_s_110_0, n1768, n213_c, ram_s_231_7, 
        n2743, n2571, n12827, ram_s_121_4, ram_s_120_4, n12830, 
        ram_s_231_6, n2742, ram_s_231_5, n2741, ram_s_231_4, n2740, 
        n2935, ram_s_255_7, n2934, ram_s_255_6, n2933, ram_s_255_5, 
        n2932, ram_s_255_4, n2931, ram_s_255_3, n2930, n2929, ram_s_255_1, 
        n2928, n2927, ram_s_254_7, n2926, ram_s_254_6, n2925, ram_s_254_5, 
        n2924, ram_s_254_4, n2923, ram_s_254_3, n2922, n2921, ram_s_254_1, 
        n2920, n2919, ram_s_253_7, n2918, ram_s_253_6, n2917, ram_s_253_5, 
        n2916, ram_s_253_4, n2915, ram_s_253_3, n2914, n2913, ram_s_253_1, 
        n2912, n2911, ram_s_252_7, n2910, ram_s_252_6, n2909, ram_s_252_5, 
        n2908, ram_s_252_4, n2907, ram_s_252_3, n2906, n2905, ram_s_252_1, 
        n2904, n2903, ram_s_251_7, n2902, n2901, ram_s_251_5, n2900, 
        n2899, ram_s_251_3, n2898, n2897, ram_s_251_1, n2896, ram_s_251_0, 
        n2895, ram_s_250_7, n2894, n2893, ram_s_250_5, n2892, n2891, 
        ram_s_250_3, n2890, n2889, ram_s_250_1, n2888, ram_s_250_0, 
        n2887, ram_s_249_7, n2886, n2885, ram_s_249_5, n2884, n2883, 
        ram_s_249_3, n2882, n2881, ram_s_249_1, n2880, ram_s_249_0, 
        n2879, ram_s_248_7, n2878, n2877, ram_s_248_5, n2876, n2875, 
        ram_s_248_3, n2874, n2873, ram_s_248_1, n2872, ram_s_248_0, 
        n2871, ram_s_247_7, n2870, ram_s_247_6, n2869, n2868, ram_s_247_4, 
        n2867, ram_s_247_3, n2866, ram_s_247_2, n2865, ram_s_247_1, 
        n2864, ram_s_247_0, n2863, ram_s_246_7, n2862, ram_s_246_6, 
        n2861, n2860, ram_s_246_4, n2859, ram_s_246_3, n2858, ram_s_246_2, 
        n2857, ram_s_246_1, n2856, ram_s_246_0, n2855, ram_s_245_7, 
        n2854, ram_s_245_6, n2853, n2852, ram_s_245_4, n2851, ram_s_245_3, 
        n2850, ram_s_245_2, n2849, ram_s_245_1, n2848, ram_s_245_0, 
        n2847, ram_s_244_7, n2846, ram_s_244_6, n2845, n2844, ram_s_244_4, 
        n2843, ram_s_244_3, n2842, ram_s_244_2, n2841, ram_s_244_1, 
        n2840, ram_s_244_0, n2839, ram_s_243_7, n2838, ram_s_243_6, 
        n2837, ram_s_243_5, n2836, ram_s_243_4, n2835, ram_s_243_3, 
        n2834, ram_s_243_2, n2833, ram_s_243_1, n2832, ram_s_243_0, 
        n2831, ram_s_242_7, n2830, ram_s_242_6, n2829, ram_s_242_5, 
        n2828, ram_s_242_4, n2827, ram_s_242_3, n2826, ram_s_242_2, 
        n2825, ram_s_242_1, n2824, ram_s_242_0, n2823, ram_s_241_7, 
        n2822, ram_s_241_6, n2821, ram_s_241_5, n2820, ram_s_241_4, 
        n2819, ram_s_241_3, n2818, ram_s_241_2, n2817, ram_s_241_1, 
        n2816, ram_s_241_0, n2815, ram_s_240_7, n2814, ram_s_240_6, 
        n2813, ram_s_240_5, n2812, ram_s_240_4, n2811, ram_s_240_3, 
        n2810, ram_s_240_2, n2809, ram_s_240_1, n2808, ram_s_240_0, 
        n2807, ram_s_239_7, n2806, ram_s_239_6, n2805, ram_s_239_5, 
        n2804, ram_s_239_4, n2803, ram_s_239_3, n2802, ram_s_239_2, 
        n2801, ram_s_239_1, n2800, ram_s_239_0, n2799, ram_s_238_7, 
        n2798, ram_s_238_6, n2797, ram_s_238_5, n2796, ram_s_238_4, 
        n2795, ram_s_238_3, n2794, ram_s_238_2, n2793, ram_s_238_1, 
        n2792, ram_s_238_0, n2739, ram_s_231_3, n2738, ram_s_231_2, 
        n2737, ram_s_231_1, n2736, ram_s_231_0, n2735, ram_s_230_7, 
        n2734, ram_s_230_6, n2733, ram_s_230_5, n2732, ram_s_230_4, 
        n2731, ram_s_230_3, n2730, ram_s_230_2, n2729, ram_s_230_1, 
        n2728, ram_s_230_0, n2727, ram_s_229_7, n2726, ram_s_229_6, 
        n2725, ram_s_229_5, n2724, ram_s_229_4, n2723, ram_s_229_3, 
        n2722, ram_s_229_2, n2721, ram_s_229_1, n2720, ram_s_229_0, 
        n2719, ram_s_228_7, n2718, ram_s_228_6, n2717, ram_s_228_5, 
        n2716, ram_s_228_4, n2715, ram_s_228_3, n2714, ram_s_228_2, 
        n2713, ram_s_228_1, n2712, ram_s_228_0, n2711, ram_s_227_7, 
        n2710, ram_s_227_6, n2709, ram_s_227_5, n2708, ram_s_227_4, 
        n2707, ram_s_227_3, n2706, ram_s_227_2, n2705, ram_s_227_1, 
        n2704, ram_s_227_0, n2703, ram_s_226_7, n2702, ram_s_226_6, 
        n2701, ram_s_226_5, n2700, ram_s_226_4, n2699, ram_s_226_3, 
        n2698, ram_s_226_2, n2697, ram_s_226_1, n2696, ram_s_226_0, 
        n2695, ram_s_225_7, n2694, ram_s_225_6, n2693, ram_s_225_5, 
        n2692, ram_s_225_4, n2691, ram_s_225_3, n2690, ram_s_225_2, 
        n2689, ram_s_225_1, n2688, ram_s_225_0, n2687, ram_s_224_7, 
        n2686, ram_s_224_6, n2685, ram_s_224_5, n2684, ram_s_224_4, 
        n2683, ram_s_224_3, n2682, ram_s_224_2, n2681, ram_s_224_1, 
        n2680, ram_s_224_0, n2679, ram_s_223_7, n2678, ram_s_223_6, 
        n2677, ram_s_223_5, n2676, ram_s_223_4, n2675, ram_s_223_3, 
        n2674, ram_s_223_2, n2673, ram_s_223_1, n2672, ram_s_223_0, 
        n2671, ram_s_222_7, n2670, ram_s_222_6, n2669, ram_s_222_5, 
        n2668, ram_s_222_4, n2667, ram_s_222_3, n2666, ram_s_222_2, 
        n2665, ram_s_222_1, n2664, ram_s_222_0, n2663, ram_s_221_7, 
        n2662, ram_s_221_6, n2661, ram_s_221_5, n2660, ram_s_221_4, 
        n2659, ram_s_221_3, n2658, ram_s_221_2, n2657, ram_s_221_1, 
        n2656, ram_s_221_0, n2655, ram_s_220_7, n2654, ram_s_220_6, 
        n2653, ram_s_220_5, n2652, ram_s_220_4, n2651, ram_s_220_3, 
        n2650, ram_s_220_2, n2649, ram_s_220_1, n2648, ram_s_220_0, 
        n2647, ram_s_219_7, n2646, ram_s_219_6, n2645, ram_s_219_5, 
        n2644, ram_s_219_4, n2643, ram_s_219_3, n2642, ram_s_219_2, 
        n2641, ram_s_219_1, n2640, ram_s_219_0, n2639, ram_s_218_7, 
        n2638, ram_s_218_6, n2637, ram_s_218_5, n2636, ram_s_218_4, 
        n2635, ram_s_218_3, n2634, ram_s_218_2, n2633, ram_s_218_1, 
        n2632, ram_s_218_0, n2631, ram_s_217_7, n2630, ram_s_217_6, 
        n2629, ram_s_217_5, n2628, ram_s_217_4, n2627, ram_s_217_3, 
        n2626, ram_s_217_2, n2625, ram_s_217_1, n2624, ram_s_217_0, 
        n2623, ram_s_216_7, n2622, ram_s_216_6, n2621, ram_s_216_5, 
        n2620, ram_s_216_4, n2619, ram_s_216_3, n2618, ram_s_216_2, 
        n2617, ram_s_216_1, n2616, ram_s_216_0, n2615, n2614, ram_s_215_6, 
        n2613, ram_s_215_5, n2612, ram_s_215_4, n2611, ram_s_215_3, 
        n2610, ram_s_215_2, n2609, ram_s_215_1, n2608, ram_s_215_0, 
        n2607, n2606, ram_s_214_6, n2605, ram_s_214_5, n2604, ram_s_214_4, 
        n2603, ram_s_214_3, n2602, ram_s_214_2, n2601, ram_s_214_1, 
        n2600, ram_s_214_0, n2599, n2598, ram_s_213_6, n2597, ram_s_213_5, 
        n2596, ram_s_213_4, n2595, ram_s_213_3, n2594, ram_s_213_2, 
        n2593, ram_s_213_1, n2592, ram_s_213_0, n2591, n2590, ram_s_212_6, 
        n2589, ram_s_212_5, n2588, ram_s_212_4, n2587, ram_s_212_3, 
        n2586, ram_s_212_2, n2585, ram_s_212_1, n2584, ram_s_212_0, 
        n2570, ram_s_210_2, n2569, ram_s_210_1, n2568, ram_s_210_0, 
        n2559, ram_s_208_7, n2558, ram_s_208_6, n2557, ram_s_208_5, 
        n2556, ram_s_208_4, n2555, n2554, ram_s_208_2, n2553, ram_s_208_1, 
        n2552, ram_s_208_0, n2549, ram_s_207_5, n2548, ram_s_207_4, 
        n2547, ram_s_207_3, n2546, ram_s_207_2, n2545, ram_s_207_1, 
        n2544, ram_s_207_0, n2543, n2542, ram_s_206_6, n2541, ram_s_206_5, 
        n2540, ram_s_206_4, n2539, ram_s_206_3, n2538, ram_s_206_2, 
        n2537, ram_s_206_1, n2536, ram_s_206_0, n2535, n2534, ram_s_205_6, 
        n2533, ram_s_205_5, n2532, ram_s_205_4, n2531, ram_s_205_3, 
        n2530, ram_s_205_2, n2529, ram_s_205_1, n2528, ram_s_205_0, 
        n2527, n2526, ram_s_204_6, n2525, ram_s_204_5, n2524, ram_s_204_4, 
        n2523, ram_s_204_3, n2522, ram_s_204_2, n2521, ram_s_204_1, 
        n2520, ram_s_204_0, n2407, n2406, ram_s_189_6, n2405, n2404, 
        ram_s_189_4, n2403, ram_s_189_3, n2402, n2401, ram_s_189_1, 
        n2400, ram_s_189_0, n2399, n2398, ram_s_188_6, n2397, n2396, 
        ram_s_188_4, n2395, ram_s_188_3, n2394, n2393, ram_s_188_1, 
        n2392, ram_s_188_0, n2391, ram_s_187_7, n2390, ram_s_187_6, 
        n2389, ram_s_187_5, n2388, ram_s_187_4, n2387, n2386, ram_s_187_2, 
        n2385, ram_s_187_1, n2384, ram_s_187_0, n2367, ram_s_184_7, 
        n2366, ram_s_184_6, n2365, ram_s_184_5, n2364, ram_s_184_4, 
        n2363, n2362, ram_s_184_2, n2361, ram_s_184_1, n2360, ram_s_184_0, 
        n2359, ram_s_183_7, n2358, ram_s_183_6, n2357, ram_s_183_5, 
        n2356, ram_s_183_4, n2355, ram_s_183_3, n2354, n2353, ram_s_183_1, 
        n2352, ram_s_183_0, n2351, ram_s_182_7, n2350, ram_s_182_6, 
        n2349, ram_s_182_5, n2348, ram_s_182_4, n2347, ram_s_182_3, 
        n2346, n2345, ram_s_182_1, n2344, ram_s_182_0, n2343, ram_s_181_7, 
        n2342, ram_s_181_6, n2341, ram_s_181_5, n2340, ram_s_181_4, 
        n2339, ram_s_181_3, n2338, n2337, ram_s_181_1, n2336, ram_s_181_0, 
        n2335, ram_s_180_7, n2334, ram_s_180_6, n2333, ram_s_180_5, 
        n2332, ram_s_180_4, n2331, ram_s_180_3, n2330, n2329, ram_s_180_1, 
        n2328, ram_s_180_0, n2327, ram_s_179_7, n2326, n2325, ram_s_179_5, 
        n2324, ram_s_179_4, n2323, ram_s_179_3, n2322, n2321, ram_s_179_1, 
        n2320, ram_s_179_0, n2319, ram_s_178_7, n2318, n2317, ram_s_178_5, 
        n2316, ram_s_178_4, n2315, ram_s_178_3, n2314, n2313, ram_s_178_1, 
        n2312, ram_s_178_0, n2311, ram_s_177_7, n2310, n2309, ram_s_177_5, 
        n2308, ram_s_177_4, n2307, ram_s_177_3, n2306, n2305, ram_s_177_1, 
        n2304, ram_s_177_0, n2303, ram_s_176_7, n2302, n2301, ram_s_176_5, 
        n2300, ram_s_176_4, n2299, ram_s_176_3, n2298, n2297, ram_s_176_1, 
        n2296, ram_s_176_0, n2287, ram_s_174_7, n2286, ram_s_174_6, 
        n2285, ram_s_174_5, n2284, ram_s_174_4, n2283, ram_s_174_3, 
        n2282, ram_s_174_2, n2281, ram_s_174_1, n2280, ram_s_174_0, 
        n2255, ram_s_170_7, n2254, ram_s_170_6, n2253, n2252, ram_s_170_4, 
        n2251, ram_s_170_3, n2250, ram_s_170_2, n2249, ram_s_170_1, 
        n2248, ram_s_170_0, n2247, ram_s_169_7, n2246, ram_s_169_6, 
        n2245, n2244, ram_s_169_4, n2243, ram_s_169_3, n2242, ram_s_169_2, 
        n2241, ram_s_169_1, n2240, ram_s_169_0, n2167, ram_s_159_7, 
        n2166, n2165, ram_s_159_5, n2164, ram_s_159_4, n2163, ram_s_159_3, 
        n2162, ram_s_159_2, n2161, n2160, ram_s_159_0, n2159, ram_s_158_7, 
        n2158, n2157, ram_s_158_5, n2156, ram_s_158_4, n2155, ram_s_158_3, 
        n2154, ram_s_158_2, n2153, n2152, ram_s_158_0, n2151, ram_s_157_7, 
        n2150, n2149, ram_s_157_5, n2148, ram_s_157_4, n2147, ram_s_157_3, 
        n2146, ram_s_157_2, n2145, n2144, ram_s_157_0, n2143, ram_s_156_7, 
        n2142, n2141, ram_s_156_5, n2140, ram_s_156_4, n2139, ram_s_156_3, 
        n2138, ram_s_156_2, n2137, n2136, ram_s_156_0, n2135, ram_s_155_7, 
        n2134, n2133, ram_s_155_5, n2132, ram_s_155_4, n2131, ram_s_155_3, 
        n2130, ram_s_155_2, n2129, ram_s_155_1, n2128, ram_s_155_0, 
        n2127, ram_s_154_7, n2126, n2125, ram_s_154_5, n2124, ram_s_154_4, 
        n2123, ram_s_154_3, n2122, ram_s_154_2, n2121, ram_s_154_1, 
        n2120, ram_s_154_0, n2119, ram_s_153_7, n2118, n2117, ram_s_153_5, 
        n2116, ram_s_153_4, n2115, ram_s_153_3, n2114, ram_s_153_2, 
        n2113, ram_s_153_1, n2112, ram_s_153_0, n2111, ram_s_152_7, 
        n2110, n2109, ram_s_152_5, n2108, ram_s_152_4, n2107, ram_s_152_3, 
        n2106, ram_s_152_2, n2105, ram_s_152_1, n2104, ram_s_152_0, 
        n2103, ram_s_151_7, n2102, ram_s_151_6, n2101, ram_s_151_5, 
        n2100, ram_s_151_4, n2099, ram_s_151_3, n2098, ram_s_151_2, 
        n2097, ram_s_151_1, n2096, ram_s_151_0, n2095, ram_s_150_7, 
        n2094, ram_s_150_6, n2093, ram_s_150_5, n2092, ram_s_150_4, 
        n2091, ram_s_150_3, n2090, ram_s_150_2, n2089, ram_s_150_1, 
        n2088, ram_s_150_0, n2087, ram_s_149_7, n2086, ram_s_149_6, 
        n2085, ram_s_149_5, n2084, ram_s_149_4, n2083, ram_s_149_3, 
        n2082, ram_s_149_2, n2081, ram_s_149_1, n2080, ram_s_149_0, 
        n2079, ram_s_148_7, n2078, ram_s_148_6, n2077, ram_s_148_5, 
        n2076, ram_s_148_4, n2075, ram_s_148_3, n2074, ram_s_148_2, 
        n2073, ram_s_148_1, n2072, ram_s_148_0, n2071, n2070, ram_s_147_6, 
        n2069, ram_s_147_5, n2068, ram_s_147_4, n2067, ram_s_147_3, 
        n2066, ram_s_147_2, n2065, ram_s_147_1, n2064, ram_s_147_0, 
        n2063, n2062, ram_s_146_6, n2061, ram_s_146_5, n2060, ram_s_146_4, 
        n2059, ram_s_146_3, n2058, ram_s_146_2, n2057, ram_s_146_1, 
        n2056, ram_s_146_0, n2055, n2054, ram_s_145_6, n2053, ram_s_145_5, 
        n2052, ram_s_145_4, n2051, ram_s_145_3, n2050, ram_s_145_2, 
        n2049, ram_s_145_1, n2048, ram_s_145_0, n2047, n2046, ram_s_144_6, 
        n2045, ram_s_144_5, n2044, ram_s_144_4, n2043, ram_s_144_3, 
        n2042, ram_s_144_2, n2041, ram_s_144_1, n2040, ram_s_144_0, 
        n2039, n2038, ram_s_143_6, n2037, n2036, ram_s_143_4, n2035, 
        n2034, ram_s_143_2, n2033, ram_s_143_1, n2032, ram_s_143_0, 
        n1999, ram_s_138_7, n1998, ram_s_138_6, n1997, ram_s_138_5, 
        n1996, ram_s_138_4, n1995, ram_s_138_3, n1994, ram_s_138_2, 
        n1993, n1992, n1991, ram_s_137_7, n1990, ram_s_137_6, n1989, 
        ram_s_137_5, n1988, ram_s_137_4, n1987, ram_s_137_3, n1986, 
        ram_s_137_2, n1985, n1984, n1911, ram_s_127_7, n1910, ram_s_127_6, 
        n1909, ram_s_127_5, n1908, ram_s_127_4, n1907, ram_s_127_3, 
        n1906, ram_s_127_2, n1905, ram_s_127_1, n1904, n1903, ram_s_126_7, 
        n1902, ram_s_126_6, n1901, ram_s_126_5, n1900, ram_s_126_4, 
        n1899, ram_s_126_3, n1898, ram_s_126_2, n1897, ram_s_126_1, 
        n1896, n1895, ram_s_125_7, n1894, ram_s_125_6, n1893, ram_s_125_5, 
        n1892, ram_s_125_4, n1891, ram_s_125_3, n1890, ram_s_125_2, 
        n1889, ram_s_125_1, n1888, n1887, ram_s_124_7, n1886, ram_s_124_6, 
        n1885, ram_s_124_5, n1884, ram_s_124_4, n1883, ram_s_124_3, 
        n1882, ram_s_124_2, n1881, ram_s_124_1, n1880, n1879, ram_s_123_7, 
        n1878, ram_s_123_6, n1877, ram_s_123_5, n1876, n1875, ram_s_123_3, 
        n1874, ram_s_123_2, n1873, ram_s_123_1, n1872, ram_s_123_0, 
        n1871, ram_s_122_7, n1870, ram_s_122_6, n1869, ram_s_122_5, 
        n1868, n1867, ram_s_122_3, n1866, ram_s_122_2, n1865, ram_s_122_1, 
        n1864, ram_s_122_0, n1863, ram_s_121_7, n1862, ram_s_121_6, 
        n1861, ram_s_121_5, n1860, n1859, ram_s_121_3, n1858, ram_s_121_2, 
        n1857, ram_s_121_1, n1856, ram_s_121_0, n1855, ram_s_120_7, 
        n1854, ram_s_120_6, n1853, ram_s_120_5, n1852, n1851, ram_s_120_3, 
        n1850, ram_s_120_2, n1849, ram_s_120_1, n1848, ram_s_120_0, 
        n1847, ram_s_119_7, n1846, ram_s_119_6, n1845, ram_s_119_5, 
        n1844, n1843, ram_s_119_3, n1842, ram_s_119_2, n1841, ram_s_119_1, 
        n1840, ram_s_119_0, n1839, ram_s_118_7, n1838, ram_s_118_6, 
        n1837, ram_s_118_5, n1836, n1835, ram_s_118_3, n1834, ram_s_118_2, 
        n1833, ram_s_118_1, n1832, ram_s_118_0, n1831, ram_s_117_7, 
        n1830, ram_s_117_6, n1829, ram_s_117_5, n1828, n1827, ram_s_117_3, 
        n1826, ram_s_117_2, n1825, ram_s_117_1, n1824, ram_s_117_0, 
        n1823, ram_s_116_7, n1822, ram_s_116_6, n1821, ram_s_116_5, 
        n1820, n1819, ram_s_116_3, n1818, ram_s_116_2, n1817, ram_s_116_1, 
        n1816, ram_s_116_0, n1767, ram_s_109_7, n1766, ram_s_109_6, 
        n1765, ram_s_109_5, n1764, ram_s_109_4, n1763, n1762, ram_s_109_2, 
        n1761, ram_s_109_1, n1760, ram_s_109_0, n1759, ram_s_108_7, 
        n1758, ram_s_108_6, n1757, ram_s_108_5, n1756, ram_s_108_4, 
        n1755, n1754, ram_s_108_2, n1753, ram_s_108_1, n1752, ram_s_108_0, 
        n1751, ram_s_107_7, n1750, ram_s_107_6, n1749, ram_s_107_5, 
        n1748, ram_s_107_4, n1747, ram_s_107_3, n1746, ram_s_107_2, 
        n1745, ram_s_107_1, n1744, ram_s_107_0, n1743, ram_s_106_7, 
        n1742, ram_s_106_6, n1741, ram_s_106_5, n1740, ram_s_106_4, 
        n1739, ram_s_106_3, n1738, ram_s_106_2, n1737, ram_s_106_1, 
        n1736, ram_s_106_0, n1735, ram_s_105_7, n1734, ram_s_105_6, 
        n1733, ram_s_105_5, n1732, ram_s_105_4, n1731, ram_s_105_3, 
        n1730, ram_s_105_2, n1729, ram_s_105_1, n1728, ram_s_105_0, 
        n1727, ram_s_104_7, n1726, ram_s_104_6, n1725, ram_s_104_5, 
        n1724, ram_s_104_4, n1723, ram_s_104_3, n1722, ram_s_104_2, 
        n1721, ram_s_104_1, n1720, ram_s_104_0, n1719, ram_s_103_7, 
        n1718, ram_s_103_6, n1717, ram_s_103_5, n1716, ram_s_103_4, 
        n1715, ram_s_103_3, n1714, ram_s_103_2, n1713, ram_s_103_1, 
        n1712, ram_s_103_0, n1711, ram_s_102_7, n1710, ram_s_102_6, 
        n1709, ram_s_102_5, n1708, ram_s_102_4, n1707, ram_s_102_3, 
        n1706, ram_s_102_2, n1705, ram_s_102_1, n1704, ram_s_102_0, 
        n1703, ram_s_101_7, n1702, ram_s_101_6, n1701, ram_s_101_5, 
        n1700, ram_s_101_4, n1699, ram_s_101_3, n1698, ram_s_101_2, 
        n1697, ram_s_101_1, n1696, ram_s_101_0, n1695, ram_s_100_7, 
        n1694, ram_s_100_6, n1693, ram_s_100_5, n1692, ram_s_100_4, 
        n1691, ram_s_100_3, n1690, ram_s_100_2, n1689, ram_s_100_1, 
        n1688, ram_s_100_0, n1687, ram_s_99_7, n1686, ram_s_99_6, 
        n1685, ram_s_99_5, n1684, ram_s_99_4, n1683, ram_s_99_3, 
        n1682, ram_s_99_2, n1681, ram_s_99_1, n1680, ram_s_99_0, 
        n1679, ram_s_98_7, n1678, ram_s_98_6, n1677, ram_s_98_5, 
        n1676, ram_s_98_4, n1675, ram_s_98_3, n1674, ram_s_98_2, 
        n1673, ram_s_98_1, n1672, ram_s_98_0, n1671, ram_s_97_7, 
        n1670, ram_s_97_6, n1669, ram_s_97_5, n1668, ram_s_97_4, 
        n1667, ram_s_97_3, n1666, ram_s_97_2, n1665, ram_s_97_1, 
        n1664, ram_s_97_0, n1663, ram_s_96_7, n1662, ram_s_96_6, 
        n1661, ram_s_96_5, n1660, ram_s_96_4, n1659, ram_s_96_3, 
        n1658, ram_s_96_2, n1657, ram_s_96_1, n1656, ram_s_96_0, 
        n1655, ram_s_95_7, n1654, n1653, n1652, ram_s_95_4, n1651, 
        ram_s_95_3, n1650, ram_s_95_2, n1649, ram_s_95_1, n1648, 
        ram_s_95_0, n1647, ram_s_94_7, n1646, n1645, n1644, ram_s_94_4, 
        n1643, ram_s_94_3, n1642, ram_s_94_2, n1641, ram_s_94_1, 
        n1640, ram_s_94_0, n1639, ram_s_93_7, n1638, n1637, n1636, 
        ram_s_93_4, n1635, ram_s_93_3, n1634, ram_s_93_2, n1633, 
        ram_s_93_1, n1632, ram_s_93_0, n1631, ram_s_92_7, n1630, 
        n1629, n1628, ram_s_92_4, n1627, ram_s_92_3, n1626, ram_s_92_2, 
        n1625, ram_s_92_1, n1624, ram_s_92_0, n1623, ram_s_91_7, 
        n1622, ram_s_91_6, n1621, ram_s_91_5, n1620, ram_s_91_4, 
        n1619, ram_s_91_3, n1618, ram_s_91_2, n1617, ram_s_91_1, 
        n1616, ram_s_91_0, n1615, ram_s_90_7, n1614, ram_s_90_6, 
        n1613, ram_s_90_5, n1612, ram_s_90_4, n1611, ram_s_90_3, 
        n1610, ram_s_90_2, n1609, ram_s_90_1, n1608, ram_s_90_0, 
        n1607, ram_s_89_7, n1606, ram_s_89_6, n1605, ram_s_89_5, 
        n1604, ram_s_89_4, n1603, ram_s_89_3, n1602, ram_s_89_2, 
        n1601, ram_s_89_1, n1600, ram_s_89_0, n1599, ram_s_88_7, 
        n1598, ram_s_88_6, n1597, ram_s_88_5, n1596, ram_s_88_4, 
        n1595, ram_s_88_3, n1594, ram_s_88_2, n1593, ram_s_88_1, 
        n1592, ram_s_88_0, n1591, n1590, ram_s_87_6, n1589, ram_s_87_5, 
        n1588, ram_s_87_4, n1587, ram_s_87_3, n1586, ram_s_87_2, 
        n1585, ram_s_87_1, n1584, ram_s_87_0, n1583, n1582, ram_s_86_6, 
        n1581, ram_s_86_5, n1580, ram_s_86_4, n1579, ram_s_86_3, 
        n1578, ram_s_86_2, n1577, ram_s_86_1, n1576, ram_s_86_0, 
        n1559, ram_s_83_7, n1558, ram_s_83_6, n1557, n1556, ram_s_83_4, 
        n1555, ram_s_83_3, n1554, ram_s_83_2, n1553, ram_s_83_1, 
        n1552, ram_s_83_0, n1551, ram_s_82_7, n1550, ram_s_82_6, 
        n1549, n1548, ram_s_82_4, n1547, ram_s_82_3, n1546, ram_s_82_2, 
        n1545, ram_s_82_1, n1544, ram_s_82_0, n1535, ram_s_80_7, 
        n1534, ram_s_80_6, n1533, n1532, ram_s_80_4, n1531, ram_s_80_3, 
        n1530, ram_s_80_2, n1529, ram_s_80_1, n1528, ram_s_80_0, 
        n1527, ram_s_79_7, n1526, ram_s_79_6, n1525, ram_s_79_5, 
        n1524, n1523, ram_s_79_3, n1522, ram_s_79_2, n1521, ram_s_79_1, 
        n1520, ram_s_79_0, n1519, ram_s_78_7, n1518, ram_s_78_6, 
        n1517, ram_s_78_5, n1516, n1515, ram_s_78_3, n1514, ram_s_78_2, 
        n1513, ram_s_78_1, n1512, ram_s_78_0, n1511, ram_s_77_7, 
        n1510, ram_s_77_6, n1509, ram_s_77_5, n1508, n1507, ram_s_77_3, 
        n1503, ram_s_76_7, n1502, ram_s_76_6, n1501, ram_s_76_5, 
        n1500, n1499, ram_s_76_3, n1498, ram_s_76_2, n1383, ram_s_61_7, 
        n1382, ram_s_61_6, n1381, ram_s_61_5, n1380, n1379, ram_s_61_3, 
        n1378, ram_s_61_2, n1377, ram_s_61_1, n1376, n1375, ram_s_60_7, 
        n1374, ram_s_60_6, n1373, ram_s_60_5, n1372, n1371, ram_s_60_3, 
        n1370, ram_s_60_2, n1369, ram_s_60_1, n1368, n1367, ram_s_59_7, 
        n1366, ram_s_59_6, n1365, n1364, ram_s_59_4, n1363, ram_s_59_3, 
        n1362, ram_s_59_2, n1361, ram_s_59_1, n1360, n1343, ram_s_56_7, 
        n1342, ram_s_56_6, n1341, n1340, ram_s_56_4, n1339, ram_s_56_3, 
        n1338, ram_s_56_2, n1337, ram_s_56_1, n1336, n1335, ram_s_55_7, 
        n1334, ram_s_55_6, n1333, ram_s_55_5, n1332, ram_s_55_4, 
        n1331, ram_s_55_3, n1330, ram_s_55_2, n1329, ram_s_55_1, 
        n1328, ram_s_55_0, n1327, ram_s_54_7, n1326, ram_s_54_6, 
        n1325, ram_s_54_5, n1324, ram_s_54_4, n1323, ram_s_54_3, 
        n1322, ram_s_54_2, n1321, ram_s_54_1, n1320, ram_s_54_0, 
        n1319, ram_s_53_7, n1318, ram_s_53_6, n1317, ram_s_53_5, 
        n1316, ram_s_53_4, n1315, ram_s_53_3, n1314, ram_s_53_2, 
        n1313, ram_s_53_1, n1312, ram_s_53_0, n1311, ram_s_52_7, 
        n1310, ram_s_52_6, n1309, ram_s_52_5, n1308, ram_s_52_4, 
        n1307, ram_s_52_3, n1306, ram_s_52_2, n1305, ram_s_52_1, 
        n1304, ram_s_52_0, n1303, ram_s_51_7, n1302, ram_s_51_6, 
        n1301, ram_s_51_5, n176_c, ram_s_20_0, n955, n1300, ram_s_51_4, 
        ram_s_20_7, n922, n1299, ram_s_51_3, ram_s_20_6, n929, n1298, 
        ram_s_51_2, ram_s_20_5, n942, n1297, ram_s_51_1, ram_s_20_4, 
        n943, n1296, ram_s_20_3, n945, n1295, ram_s_50_7, ram_s_20_2, 
        n947, n1294, ram_s_50_6, ram_s_20_1, n954, n1293, ram_s_50_5, 
        n172, ram_s_18_2, n1024, n1292, ram_s_50_4, ram_s_18_6, 
        n1020, n1291, ram_s_50_3, ram_s_18_5, n1021, n1290, ram_s_50_2, 
        ram_s_18_4, n1022, n1289, ram_s_50_1, ram_s_18_3, n1023, 
        n1288, ram_s_18_7, n1019, n1287, ram_s_49_7, ram_s_18_1, 
        n919, n1286, ram_s_49_6, n921, n1285, ram_s_49_5, ram_s_19_2, 
        n1057, n1284, ram_s_49_4, ram_s_19_5, n1027, n1283, ram_s_49_3, 
        ram_s_19_4, n1028, n1282, ram_s_49_2, ram_s_19_3, n1050, 
        n1281, ram_s_49_1, ram_s_19_1, n914, n1280, n1018, n1279, 
        ram_s_48_7, ram_s_19_7, n1025, n1278, ram_s_48_6, ram_s_19_6, 
        n1026, n1277, ram_s_48_5, n168, n1059, n1276, ram_s_48_4, 
        ram_s_16_7, n951, n1275, ram_s_48_3, ram_s_16_6, n953, n1274, 
        ram_s_48_2, ram_s_16_5, n1048, n1273, ram_s_48_1, ram_s_16_4, 
        n1053, n1272, ram_s_16_3, n1054, ram_s_16_2, n1055, ram_s_16_1, 
        n1058, n166, ram_s_15_7, n1060, ram_s_15_4, n900, ram_s_15_3, 
        n902, ram_s_15_2, n903, ram_s_15_1, n913, ram_s_15_0, n956, 
        n1263, ram_s_46_7, n1049, n1262, ram_s_46_6, n1052, n1261, 
        ram_s_46_5, n180, ram_s_22_7, n1071, n1260, ram_s_46_4, 
        ram_s_22_6, n1070, n1259, ram_s_46_3, ram_s_22_5, n1069, 
        n1258, ram_s_22_4, n1068, n1257, ram_s_46_1, ram_s_22_3, 
        n1067, n1256, ram_s_46_0, ram_s_22_2, n1066, ram_s_22_1, 
        n1065, ram_s_22_0, n1064, n182_c, ram_s_23_7, n1079, ram_s_23_6, 
        n1078, ram_s_23_5, n1077, ram_s_23_4, n1076, ram_s_23_3, 
        n1075, ram_s_23_2, n1074, ram_s_23_1, n1073, ram_s_23_0, 
        n1072, n184_c, ram_s_24_7, n1087, ram_s_24_6, n1086, ram_s_24_5, 
        n1085, ram_s_24_4, n1084, ram_s_24_3, n1083, ram_s_24_2, 
        n1082, ram_s_24_1, n1081, ram_s_24_0, n1080, n186_c, ram_s_25_7, 
        n1095, ram_s_25_6, n1094, ram_s_25_5, n1093, ram_s_25_4, 
        n1092, ram_s_25_3, n1091, ram_s_25_2, n1090, n1231, ram_s_25_1, 
        n1089, n1230, ram_s_42_6, ram_s_25_0, n1088, n1229, ram_s_42_5, 
        n188_c, ram_s_26_7, n1103, n1228, ram_s_42_4, ram_s_26_6, 
        n1102, n1227, ram_s_42_3, ram_s_26_5, n1101, n1226, ram_s_26_4, 
        n1100, n1225, ram_s_26_3, n1099, n1224, ram_s_42_0, ram_s_26_2, 
        n1098, n1223, ram_s_26_1, n1097, n1222, ram_s_41_6, ram_s_26_0, 
        n1096, n1221, ram_s_41_5, n190_c, ram_s_27_7, n1111, n1220, 
        ram_s_41_4, ram_s_27_6, n1110, n1219, ram_s_41_3, ram_s_27_5, 
        n1109, n1218, ram_s_27_4, n1108, n1217, ram_s_27_3, n1107, 
        n1216, ram_s_41_0, ram_s_27_2, n1106, ram_s_27_1, n1105, 
        ram_s_27_0, n1104, n192_c, ram_s_28_7, n1119, ram_s_28_6, 
        n1118, n1117, ram_s_28_4, n1116, ram_s_28_3, n1115, ram_s_28_2, 
        n1114, n1113, ram_s_28_0, n1112, n194_c, ram_s_29_7, n1127, 
        ram_s_29_6, n1126, n1125, ram_s_29_4, n1124, ram_s_29_3, 
        n1123, ram_s_29_2, n1122, n1121, ram_s_29_0, n1120, n196, 
        ram_s_30_7, n1135, ram_s_30_6, n1134, n1133, ram_s_30_4, 
        n1132, ram_s_30_3, n1131, ram_s_30_2, n1130, n1129, ram_s_30_0, 
        n1128, n198, ram_s_31_7, n1143, ram_s_31_6, n1142, n1141, 
        ram_s_31_4, n1140, ram_s_31_3, n1139, ram_s_31_2, n1138, 
        n1137, ram_s_31_0, n1136, n218_c, n220_c, n228, n232, 
        n234, n236, n238, n240, n242, n244_c, n246_c, n248, 
        n254_c, n256_c, n258, n1063, ram_s_21_7, n1062, ram_s_21_6, 
        n163, n1061, ram_s_21_5, n1056, ram_s_21_4, n1039, ram_s_17_6, 
        n94_c, n92_c, n90_c, n88, n86_c, n84_c, n82_c, n80, 
        n78, n76, n74, n72_c, n133, n131, n1000, ram_s_9_3, 
        n999, ram_s_9_0, n991, ram_s_9_4, n990, ram_s_9_1, n123_c, 
        n121_c, n982, ram_s_9_5, n981, n949, ram_s_10_5, n948, 
        n928, ram_s_9_7, n101, n9375, n9376, n11465, n9352, n9351, 
        n11468, n10104, n10105, n11459, n10102, n10101, n11462, 
        n11453, n9306, n9307, n11447, n9292, n9291, n11450, n10439, 
        n10475, n11441, n10388, n11444, n11429, n11432, n11423, 
        n11426, n10613, n10631, n11417, n10601, n10580, n11420, 
        n8957, n8966, n11411, n8933, n8921, n11414, n11405, n11408, 
        n10319, n10352, n11399, n10283, n10247, n11402, n11393, 
        n11396, n11387, n11390, n11381, n11384, n9467, n11375, 
        n11366, n11330, n10562, n11369, n11372, n11363, n9639, 
        n9640, n11357, n9622, n9621, n11360, n11351, n11354, n9441, 
        n9442, n11333, n9424, n9423, n11336, n11327, n10068, n10069, 
        n11321, n10060, n10059, n11324, n11309, n11312, n11297, 
        n11291, n11294, n11285, n97_c, n11279, n11282, n11267, 
        n11270, n9234, n9235, n11255, n9217, n9216, n11258, n11249, 
        n9110, n9122, n11243, n9107, n9098, n11246, n10592, n10628, 
        n11237, n10529, n11240, n95_c, n93_c, n211, n71_adj_842, 
        n199_adj_843, n9629, n12311, n9557, n9491, n12314, n9650, 
        n11555, n9605, n9584, n11558, n12083, n12086, n12305, 
        n12308, n73, n201, n75, n203, n87, n85_adj_845, n77, 
        n205, n83, n81, n79, n207, n209, n156, n920, ram_s_17_7, 
        n915, ram_s_21_0, ram_s_10_7, n910, n11177, n27, n11180, 
        n11, n15, n16, n249_c, n251_c, n259, n21, n37, n261, 
        n10250, n8813, n11171, n43, n8798, n8855, n11174, n197, 
        n14480, n11810, n14198, n19, n35, n195_adj_858, n18, n25, 
        n154, n193_adj_859, n65_adj_860, n167, n178, n191_adj_861, 
        n63_adj_862, n12821, n10088, n170, n98, n22, n100, n96_adj_864, 
        ram_s_21_2, n905, ram_s_21_1, n912, n49, n17, n41, n257_adj_873, 
        n255_adj_874, n253_adj_875, n61_adj_876, n187_adj_877, n185_adj_878, 
        n247, n55_adj_879, n245_adj_880, n53, n243_adj_881, n51, 
        n241, n239, n189_adj_882, n47, n20, n39, n12809, n12812, 
        n10640, n10664, n12803, n10595, n10574, n12806, n12797, 
        n12800, n12791, n9710, n12785, n10826, n12773, n12776, 
        n12767, n9368, n12761, n9074, n12755, n12758, n12749, 
        n12299, n12752, n12302, n183_adj_883, n10676, n10679, n12743, 
        n10667, n10658, n10829, n12737, n12740, n12731, n9719, 
        n12293, n10412, n12077, n10394, n10370, n12080, n11696, 
        n9119, n9131, n11873, n9101, n11876, n11543, n9227, n9251, 
        n12071, n9182, n9161, n12074, n11546, n11687, n11867, 
        n11540, n11060, n11690, n11870, n12065, n9077, n11681, 
        n12059, n11684, n9728, n9737, n11537, n12062, n14450, 
        n14348, n12287, n12290, n12053, n9905, n9917, n11855, 
        n9899, n9884, n11054, n12719, n10065, n10066, n11849, 
        n12281, n12056, n12284, n10048, n10047, n11852, n11675, 
        n9278, n9941, n12275, n12047, n12050, n8825, n10646, n12278, 
        n12269, n12263, n12722, n12713, n12716, n12707, n9564, 
        n9565, n12701, n9547, n9546, n12695, n12380, n12242, n12689, 
        n12440, n12626, n12692, n12266, n12041, n11669, n11672, 
        n14090, n14006, n12044, n9959, n9980, n12677, n11837, 
        n9512, n9536, n11663, n12035, n11531, n12257, n9461, n9440, 
        n11666, n12038, n9923, n9887, n12680, n12218, n12014, 
        n12674, n12578, n8930, n8939, n12671, n8927, n12665, n12659, 
        n9594, n9595, n12653, n9586, n9585, n10712, n10715, n12647, 
        n10703, n10694, n10838, n12641, n12635, n12638, n12629, 
        n12632, n12029, n11534, n12623, n12023, n12251, n9944, 
        n9953, n11819, n9929, n9920, n11072, n10481, n12617, n12620, 
        n12017, n12611, n12605, n12608, n11639, n11642, n10457, 
        n10445, n12020, n12599, n10844, n12593, n12596, n9620, 
        n9632, n12587, n9614, n9599, n12590, n12581, n8963, n8975, 
        n12575, n8960, n8951, n12569, n10745, n10757, n12563, 
        n10739, n10721, n10847, n12245, n12248, n11633, n11636, 
        n12239, n8945, n8969, n12233, n9032, n12011, n11954, n12236, 
        n9029, n9020, n10340, n10358, n12227, n10322, n10304, 
        n12230, n9188, n9200, n11813, n11627, n12005, n9167, n9152, 
        n11816, n12008, n11786, n8935, n11807, n12221, n8917, 
        n11780, n11999, n9323, n9302, n12002, n10941, n10942, 
        n11801, n10906, n10905, n11804, n8903, n11993, n10881, 
        n11795, n10870, n10869, n11798, n11996, n9002, n9011, 
        n12215, n12557, n12560, n12551, n12554, n9714, n9715, 
        n12539, n9694, n9693, n12542, n12533, n12536, n12494, 
        n12527, n10052, n10016, n12530, n10775, n10799, n12521, 
        n10730, n10709, n12524, n8999, n8981, n11621, n12515, 
        n12518, n12509, n12497, n10815, n11789, n10786, n10785, 
        n11792, n12209, n11960, n12212, n10812, n11783, n11624, 
        n11525, n10801, n10800, n11981, n10746, n10747, n11777, 
        n10723, n10722, n11984, n11615, n11618, n10268, n11528, 
        n11771, n11609, n11975, n9272, n9206, n12500, n12491, 
        n181, n12485, n12488, n12479, n10781, n10790, n12473, 
        n13205, n13211, n13214, n10769, n10760, n10856, n12461, 
        n12464, n12164, n12455, n12422, n12458, n12449, n10793, 
        n10859, n12443, n12446, n12437, n10691, n10700, n11969, 
        n12191, n9981, n9982, n12185, n10670, n10655, n11972, 
        n9913, n9912, n12179, n12182, n12173, n12176, n12167, 
        n12170, n12161, n11963, n11765, n11768, n11612, n12155, 
        n11957, n9987, n9988, n12425, n9973, n9972, n12428, n12419, 
        n12413, n12416, n10331, n12407, n9893, n9608, n10013, 
        n10037, n12401, n9998, n9977, n12404, n12395, n12398, 
        n12158, n11951, n12143, n11603, n11753, n11597, n10718, 
        n10751, n11591, n10682, n10661, n11594, n12383, n12377, 
        n13229, n13232, n13235, n13241, n13247, n13250, n13253, 
        n9454, n9453, n13256, n9480, n9481, n13259, n13277, n13283, 
        n13286, n13289, n13295, n13298, n13301, n10577, n13307, 
        n13313, n13316, n13319, n13322, n13325, n13328, n13331, 
        n13337, n13343, n13346, n13349, n13355, n13361, n13367, 
        n13370, n13373, n13376, n13379, n13382, n13385, n13388, 
        n13391, n13397, n13403, n9509, n9479, n13406, n9545, n9581, 
        n13409, n13415, n9932, n9911, n9950, n9971, n13421, n13424, 
        n13427, n13433, n13439, n13445, n13448, n13451, n13454, 
        n13457, n8942, n8978, n13463, n13466, n13469, n13475, 
        n13478, n13481, n13487, n13493, n13499, n13511, n13517, 
        n13520, n13529, n13532, n9437, n13535, n13538, n13541, 
        n13547, n13550, n13553, n10706, n10697, n10727, n10742, 
        n13559, n10009, n10008, n13562, n10017, n10018, n13571, 
        n13577, n13580, n13583, n13589, n13592, n13595, n13601, 
        n9866, n9836, n9878, n9902, n13607, n13610, n13613, n13619, 
        n13622, n13625, n10385, n10367, n10391, n13631, n13637, 
        n13640, n13643, n13646, n13649, n13655, n13661, n13667, 
        n13673, n10619, n10685, n13679, n13682, n13685, n13691, 
        n13697, n10346, n10337, n10349, n10361, n13709, n8804, 
        n13715, n10637, n10616, n10652, n10673, n13727, n10313, 
        n10301, n10316, n10325, n13733, n13757, n13760, n13763, 
        n13766, n13769, n13775, n13778, n13781, n9806, n9827, 
        n13787, n10583, n10607, n13793, n13799, n13802, n13805, 
        n13808, n13811, n9133, n9132, n13814, n9147, n9148, n13817, 
        n9493, n9492, n13820, n9504, n9505, n13823, n13826, n13829, 
        n9124, n9123, n9156, n9157, n13841, n10271, n10256, n10277, 
        n10295, n13847, n13853, n13859, n13865, n9202, n9201, 
        n13868, n9213, n9214, n13871, n13877, n13883, n10286, 
        n13889, n13895, n10229, n10241, n10253, n13901, n13907, 
        n13913, n13916, n13919, n13925, n13928, n13931, n13934, 
        n13937, n13940, n8848, n13943, n13946, n13949, n13955, 
        n13958, n13961, n13964, n13967, n13973, n13976, n13979, 
        n13985, n13991, n13997, n14000, n14003, n14009, n14012, 
        n14021, n14027, n14030, n14033, n14039, n9487, n9486, 
        n14042, n9498, n9499, n14045, n14051, n14057, n14063, 
        n14066, n14075, n14081, n14084, n14087, n14093, n14099, 
        n14102, n14105, n14111, n14114, n14117, n14123, n14126, 
        n14129, n179, n14141, n14147, n14150, n14153, n14156, 
        n14159, n14165, n14168, n14171, n14174, n14177, n14183, 
        n14186, n14189, n14195, n8953, n8970, n8971, n14201, n14207, 
        n14213, n14216, n14219, n14225, n9842, n14231, n14237, 
        n14243, n14249, n14255, n14261, n14264, n14267, n9860, 
        n9833, n14270, n9875, n9896, n14273, n14276, n14279, n14285, 
        n14288, n14291, n10598, n9041, n14297, n14303, n14306, 
        n14309, n14312, n14315, n14321, n14327, n14333, n14339, 
        n9803, n9821, n14345, n14351, n14354, n14357, n14363, 
        n14369, n14381, n14384, n14387, n14393, n14399, n14405, 
        n14411, n14414, n14417, n14423, n14429, n14432, n14435, 
        n9140, n9515, n14447, n14453, n14456, n14459, n14465, 
        n14471, n14477, n9502, n9501, n9517, n14483, n14486, n14489, 
        n14495, n14501, n14507, n9472, n9475, n14513, n14519, 
        n14525, n14528, n14531, n14537, n14543, n14549, n14552, 
        n14555, n14561, n14567, n14573, n14585, n14591, n14594, 
        n14597, n9428, n9449, n9458, n14603, n14609, n14612, n14615, 
        n14621, n14624, n14627, n14633, n14639, n14645, n14657, 
        n14663, n14669, n14675, n14681, n14684, n14687, n14690, 
        n9847, n14693, n9430, n9433, n14699, n14702, n14705, n14708, 
        n14711, n14717, n10232, n10259, n10274, n14723, n14729, 
        n14735, n14741, n14747, n14753, n14759, n14765, n14777, 
        n14789, n14795, n14801, n14804, n14807, n14813, n14819, 
        n14825, n14831, n14837, n14843, n14849, n14855, n14861, 
        n14867, n14873, n14879, n9824, n9812, n9830, n9851, n14885, 
        n14891, n14894, n14897, n14909, n14915, n14921, n14927, 
        n14930, n14933, n8843, n14939, n14945, n14951, n14957, 
        n14963, n14975, n14981, n14987, n14993, n14999, n15005, 
        n15011, n15017, n15029, n15035, n15041, n15047, n15053, 
        n15059, n15062, n15065, n15071, n15077, n15083, n15089, 
        n15095, n15101, n15107, n15113, n15119, n15125, n15128, 
        n15131, n15137, n15143, n9104, n9113, n15149, n15155, 
        n15161, n10238, n15167, n15173, n15179, n15185, n15191, 
        n15197, n15203, n15209, n15212, n15215, n15221, n15227, 
        n15233, n15245, n15251, n15257, n15263, n15269, n15275, 
        n15281, n15287, n15293, n15299, n15305, n15311, n15317, 
        n8812, n9277, n8824, n9931, n8941, n8977, n9865, n9835, 
        n9040, n8842;
    
    SB_LUT4 port_id_0__bdd_4_lut_11798 (.I0(port_id[0]), .I1(ram_s_70_3), 
            .I2(ram_s_71_3), .I3(port_id[1]), .O(n13199));
    defparam port_id_0__bdd_4_lut_11798.LUT_INIT = 16'he4aa;
    SB_LUT4 n13199_bdd_4_lut (.I0(n13199), .I1(ram_s_69_3), .I2(ram_s_68_3), 
            .I3(port_id[1]), .O(n9038));
    defparam n13199_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11793 (.I0(port_id[0]), .I1(ram_s_154_6), 
            .I2(ram_s_155_6), .I3(port_id[1]), .O(n13193));
    defparam port_id_0__bdd_4_lut_11793.LUT_INIT = 16'he4aa;
    SB_LUT4 n13193_bdd_4_lut (.I0(n13193), .I1(ram_s_153_6), .I2(ram_s_152_6), 
            .I3(port_id[1]), .O(n13196));
    defparam n13193_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11788 (.I0(port_id[0]), .I1(ram_s_254_0), 
            .I2(ram_s_255_0), .I3(port_id[1]), .O(n13187));
    defparam port_id_0__bdd_4_lut_11788.LUT_INIT = 16'he4aa;
    SB_LUT4 n13187_bdd_4_lut (.I0(n13187), .I1(ram_s_253_0), .I2(ram_s_252_0), 
            .I3(port_id[1]), .O(n13190));
    defparam n13187_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1327_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_85_7), .O(n1575));   // src/ram.vhd(68[19:45])
    defparam i1327_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1567_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_115_7), .O(n1815));   // src/ram.vhd(68[19:45])
    defparam i1567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1326_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_85_6), .O(n1574));   // src/ram.vhd(68[19:45])
    defparam i1326_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1566_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_115_6), .O(n1814));   // src/ram.vhd(68[19:45])
    defparam i1566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1565_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_115_5), .O(n1813));   // src/ram.vhd(68[19:45])
    defparam i1565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1564_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_115_4), .O(n1812));   // src/ram.vhd(68[19:45])
    defparam i1564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1258_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_77_2), .O(n1506));   // src/ram.vhd(68[19:45])
    defparam i1258_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11783 (.I0(port_id[0]), .I1(ram_s_34_7), 
            .I2(ram_s_35_7), .I3(port_id[1]), .O(n13181));
    defparam port_id_0__bdd_4_lut_11783.LUT_INIT = 16'he4aa;
    SB_LUT4 n13181_bdd_4_lut (.I0(n13181), .I1(ram_s_33_7), .I2(ram_s_32_7), 
            .I3(port_id[1]), .O(n13184));
    defparam n13181_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1249_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_76_1), .O(n1497));   // src/ram.vhd(68[19:45])
    defparam i1249_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11778 (.I0(port_id[0]), .I1(ram_s_10_6), 
            .I2(ram_s_11_6), .I3(port_id[1]), .O(n13175));
    defparam port_id_0__bdd_4_lut_11778.LUT_INIT = 16'he4aa;
    SB_LUT4 n13175_bdd_4_lut (.I0(n13175), .I1(ram_s_9_6), .I2(ram_s_8_6), 
            .I3(port_id[1]), .O(n9044));
    defparam n13175_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1325_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_85_5), .O(n1573));   // src/ram.vhd(68[19:45])
    defparam i1325_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1563_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_115_3), .O(n1811));   // src/ram.vhd(68[19:45])
    defparam i1563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_5__bdd_4_lut_12622 (.I0(port_id[5]), .I1(n9495), .I2(n9496), 
            .I3(port_id[6]), .O(n13169));
    defparam port_id_5__bdd_4_lut_12622.LUT_INIT = 16'he4aa;
    SB_LUT4 n13169_bdd_4_lut (.I0(n13169), .I1(n9484), .I2(n9483), .I3(port_id[6]), 
            .O(n13172));
    defparam n13169_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11773 (.I0(port_id[0]), .I1(ram_s_250_2), 
            .I2(ram_s_251_2), .I3(port_id[1]), .O(n13163));
    defparam port_id_0__bdd_4_lut_11773.LUT_INIT = 16'he4aa;
    SB_LUT4 i1562_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_115_2), .O(n1810));   // src/ram.vhd(68[19:45])
    defparam i1562_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13163_bdd_4_lut (.I0(n13163), .I1(ram_s_249_2), .I2(ram_s_248_2), 
            .I3(port_id[1]), .O(n13166));
    defparam n13163_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1324_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_85_4), .O(n1572));   // src/ram.vhd(68[19:45])
    defparam i1324_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11763 (.I0(port_id[0]), .I1(ram_s_126_0), 
            .I2(ram_s_127_0), .I3(port_id[1]), .O(n13157));
    defparam port_id_0__bdd_4_lut_11763.LUT_INIT = 16'he4aa;
    SB_LUT4 i1561_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_115_1), .O(n1809));   // src/ram.vhd(68[19:45])
    defparam i1561_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13157_bdd_4_lut (.I0(n13157), .I1(ram_s_125_0), .I2(ram_s_124_0), 
            .I3(port_id[1]), .O(n9047));
    defparam n13157_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut_12407 (.I0(port_id[3]), .I1(n13004), .I2(n9451), 
            .I3(port_id[4]), .O(n13151));
    defparam port_id_3__bdd_4_lut_12407.LUT_INIT = 16'he4aa;
    SB_LUT4 n13151_bdd_4_lut (.I0(n13151), .I1(n9445), .I2(n12992), .I3(port_id[4]), 
            .O(n13154));
    defparam n13151_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_6__bdd_4_lut_12008 (.I0(port_id[6]), .I1(n10025), .I2(n10043), 
            .I3(port_id[7]), .O(n13145));
    defparam port_id_6__bdd_4_lut_12008.LUT_INIT = 16'he4aa;
    SB_LUT4 n13145_bdd_4_lut (.I0(n13145), .I1(n10004), .I2(n9995), .I3(port_id[7]), 
            .O(spm_ram_data[2]));
    defparam n13145_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11758 (.I0(port_id[0]), .I1(ram_s_62_4), 
            .I2(ram_s_63_4), .I3(port_id[1]), .O(n13139));
    defparam port_id_0__bdd_4_lut_11758.LUT_INIT = 16'he4aa;
    SB_LUT4 n13139_bdd_4_lut (.I0(n13139), .I1(ram_s_61_4), .I2(ram_s_60_4), 
            .I3(port_id[1]), .O(n9671));
    defparam n13139_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11743 (.I0(port_id[0]), .I1(ram_s_2_7), 
            .I2(ram_s_3_7), .I3(port_id[1]), .O(n13133));
    defparam port_id_0__bdd_4_lut_11743.LUT_INIT = 16'he4aa;
    SB_LUT4 n13133_bdd_4_lut (.I0(n13133), .I1(ram_s_1_7), .I2(ram_s_0_7), 
            .I3(port_id[1]), .O(n13136));
    defparam n13133_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11738 (.I0(port_id[0]), .I1(ram_s_66_4), 
            .I2(ram_s_67_4), .I3(port_id[1]), .O(n13127));
    defparam port_id_0__bdd_4_lut_11738.LUT_INIT = 16'he4aa;
    SB_LUT4 n13127_bdd_4_lut (.I0(n13127), .I1(ram_s_65_4), .I2(ram_s_64_4), 
            .I3(port_id[1]), .O(n9674));
    defparam n13127_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11878 (.I0(port_id[2]), .I1(n12260), .I2(n12194), 
            .I3(port_id[3]), .O(n13121));
    defparam port_id_2__bdd_4_lut_11878.LUT_INIT = 16'he4aa;
    SB_LUT4 n13121_bdd_4_lut (.I0(n13121), .I1(n12272), .I2(n12356), .I3(port_id[3]), 
            .O(n13124));
    defparam n13121_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1560_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_115_0), .O(n1808));   // src/ram.vhd(68[19:45])
    defparam i1560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11733 (.I0(port_id[0]), .I1(ram_s_254_2), 
            .I2(ram_s_255_2), .I3(port_id[1]), .O(n13115));
    defparam port_id_0__bdd_4_lut_11733.LUT_INIT = 16'he4aa;
    SB_LUT4 n13115_bdd_4_lut (.I0(n13115), .I1(ram_s_253_2), .I2(ram_s_252_2), 
            .I3(port_id[1]), .O(n13118));
    defparam n13115_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2543_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_237_7), .O(n2791));   // src/ram.vhd(68[19:45])
    defparam i2543_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_2__bdd_4_lut_11728 (.I0(port_id[2]), .I1(n10604), .I2(n10610), 
            .I3(port_id[3]), .O(n13109));
    defparam port_id_2__bdd_4_lut_11728.LUT_INIT = 16'he4aa;
    SB_LUT4 n13109_bdd_4_lut (.I0(n13109), .I1(n10589), .I2(n10586), .I3(port_id[3]), 
            .O(n10805));
    defparam n13109_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11723 (.I0(port_id[0]), .I1(ram_s_246_5), 
            .I2(ram_s_247_5), .I3(port_id[1]), .O(n13103));
    defparam port_id_0__bdd_4_lut_11723.LUT_INIT = 16'he4aa;
    SB_LUT4 n13103_bdd_4_lut (.I0(n13103), .I1(ram_s_245_5), .I2(ram_s_244_5), 
            .I3(port_id[1]), .O(n10418));
    defparam n13103_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11713 (.I0(port_id[0]), .I1(ram_s_142_3), 
            .I2(ram_s_143_3), .I3(port_id[1]), .O(n13097));
    defparam port_id_0__bdd_4_lut_11713.LUT_INIT = 16'he4aa;
    SB_LUT4 n13097_bdd_4_lut (.I0(n13097), .I1(ram_s_141_3), .I2(ram_s_140_3), 
            .I3(port_id[1]), .O(n9680));
    defparam n13097_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2542_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_237_6), .O(n2790));   // src/ram.vhd(68[19:45])
    defparam i2542_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11708 (.I0(port_id[0]), .I1(ram_s_158_6), 
            .I2(ram_s_159_6), .I3(port_id[1]), .O(n13091));
    defparam port_id_0__bdd_4_lut_11708.LUT_INIT = 16'he4aa;
    SB_LUT4 n13091_bdd_4_lut (.I0(n13091), .I1(ram_s_157_6), .I2(ram_s_156_6), 
            .I3(port_id[1]), .O(n13094));
    defparam n13091_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2541_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_237_5), .O(n2789));   // src/ram.vhd(68[19:45])
    defparam i2541_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2540_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_237_4), .O(n2788));   // src/ram.vhd(68[19:45])
    defparam i2540_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11703 (.I0(port_id[0]), .I1(ram_s_178_2), 
            .I2(ram_s_179_2), .I3(port_id[1]), .O(n13085));
    defparam port_id_0__bdd_4_lut_11703.LUT_INIT = 16'he4aa;
    SB_LUT4 n13085_bdd_4_lut (.I0(n13085), .I1(ram_s_177_2), .I2(ram_s_176_2), 
            .I3(port_id[1]), .O(n13088));
    defparam n13085_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11838 (.I0(port_id[1]), .I1(n9336), .I2(n9337), 
            .I3(port_id[2]), .O(n13079));
    defparam port_id_1__bdd_4_lut_11838.LUT_INIT = 16'he4aa;
    SB_LUT4 i2539_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_237_3), .O(n2787));   // src/ram.vhd(68[19:45])
    defparam i2539_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13079_bdd_4_lut (.I0(n13079), .I1(n9328), .I2(n9327), .I3(port_id[2]), 
            .O(n13082));
    defparam n13079_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2538_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_237_2), .O(n2786));   // src/ram.vhd(68[19:45])
    defparam i2538_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i260_261 (.Q(ram_s_10_2), .C(CLK_3P3_MHZ_c), .D(n898));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1323_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_85_3), .O(n1571));   // src/ram.vhd(68[19:45])
    defparam i1323_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10175 (.I0(port_id[0]), .I1(ram_s_210_3), 
            .I2(ram_s_211_3), .I3(port_id[1]), .O(n11225));
    defparam port_id_0__bdd_4_lut_10175.LUT_INIT = 16'he4aa;
    SB_LUT4 i2537_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_237_1), .O(n2785));   // src/ram.vhd(68[19:45])
    defparam i2537_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11225_bdd_4_lut (.I0(n11225), .I1(ram_s_209_3), .I2(ram_s_208_3), 
            .I3(port_id[1]), .O(n11228));
    defparam n11225_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2536_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_237_0), .O(n2784));   // src/ram.vhd(68[19:45])
    defparam i2536_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1322_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_85_2), .O(n1570));   // src/ram.vhd(68[19:45])
    defparam i1322_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11698 (.I0(port_id[0]), .I1(ram_s_130_0), 
            .I2(ram_s_131_0), .I3(port_id[1]), .O(n13073));
    defparam port_id_0__bdd_4_lut_11698.LUT_INIT = 16'he4aa;
    SB_LUT4 i1321_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_85_1), .O(n1569));   // src/ram.vhd(68[19:45])
    defparam i1321_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1559_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_114_7), .O(n1807));   // src/ram.vhd(68[19:45])
    defparam i1559_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1558_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_114_6), .O(n1806));   // src/ram.vhd(68[19:45])
    defparam i1558_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13073_bdd_4_lut (.I0(n13073), .I1(ram_s_129_0), .I2(ram_s_128_0), 
            .I3(port_id[1]), .O(n9053));
    defparam n13073_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1557_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_114_5), .O(n1805));   // src/ram.vhd(68[19:45])
    defparam i1557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1556_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_114_4), .O(n1804));   // src/ram.vhd(68[19:45])
    defparam i1556_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11688 (.I0(port_id[0]), .I1(ram_s_70_4), 
            .I2(ram_s_71_4), .I3(port_id[1]), .O(n13067));
    defparam port_id_0__bdd_4_lut_11688.LUT_INIT = 16'he4aa;
    SB_LUT4 i1555_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_114_3), .O(n1803));   // src/ram.vhd(68[19:45])
    defparam i1555_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10915 (.I0(port_id[0]), .I1(ram_s_30_1), 
            .I2(ram_s_31_1), .I3(port_id[1]), .O(n12137));
    defparam port_id_0__bdd_4_lut_10915.LUT_INIT = 16'he4aa;
    SB_LUT4 n13067_bdd_4_lut (.I0(n13067), .I1(ram_s_69_4), .I2(ram_s_68_4), 
            .I3(port_id[1]), .O(n9686));
    defparam n13067_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12137_bdd_4_lut (.I0(n12137), .I1(ram_s_29_1), .I2(ram_s_28_1), 
            .I3(port_id[1]), .O(n12140));
    defparam n12137_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11683 (.I0(port_id[0]), .I1(ram_s_170_5), 
            .I2(ram_s_171_5), .I3(port_id[1]), .O(n13061));
    defparam port_id_0__bdd_4_lut_11683.LUT_INIT = 16'he4aa;
    SB_LUT4 n13061_bdd_4_lut (.I0(n13061), .I1(ram_s_169_5), .I2(ram_s_168_5), 
            .I3(port_id[1]), .O(n9347));
    defparam n13061_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11693 (.I0(port_id[1]), .I1(n9312), .I2(n9313), 
            .I3(port_id[2]), .O(n13055));
    defparam port_id_1__bdd_4_lut_11693.LUT_INIT = 16'he4aa;
    SB_LUT4 n13055_bdd_4_lut (.I0(n13055), .I1(n9304), .I2(n9303), .I3(port_id[2]), 
            .O(n13058));
    defparam n13055_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11678 (.I0(port_id[0]), .I1(ram_s_14_6), 
            .I2(ram_s_15_6), .I3(port_id[1]), .O(n13049));
    defparam port_id_0__bdd_4_lut_11678.LUT_INIT = 16'he4aa;
    SB_LUT4 n13049_bdd_4_lut (.I0(n13049), .I1(ram_s_13_6), .I2(ram_s_12_6), 
            .I3(port_id[1]), .O(n9056));
    defparam n13049_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11673 (.I0(port_id[1]), .I1(n9282), .I2(n9283), 
            .I3(port_id[2]), .O(n13043));
    defparam port_id_1__bdd_4_lut_11673.LUT_INIT = 16'he4aa;
    SB_LUT4 n13043_bdd_4_lut (.I0(n13043), .I1(n9262), .I2(n9261), .I3(port_id[2]), 
            .O(n13046));
    defparam n13043_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1554_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_114_2), .O(n1802));   // src/ram.vhd(68[19:45])
    defparam i1554_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1553_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_114_1), .O(n1801));   // src/ram.vhd(68[19:45])
    defparam i1553_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10156 (.I0(port_id[0]), .I1(ram_s_202_1), 
            .I2(ram_s_203_1), .I3(port_id[1]), .O(n11219));
    defparam port_id_0__bdd_4_lut_10156.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11110 (.I0(port_id[0]), .I1(ram_s_6_5), 
            .I2(ram_s_7_5), .I3(port_id[1]), .O(n12359));
    defparam port_id_0__bdd_4_lut_11110.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10755 (.I0(port_id[0]), .I1(ram_s_14_5), 
            .I2(ram_s_15_5), .I3(port_id[1]), .O(n11939));
    defparam port_id_0__bdd_4_lut_10755.LUT_INIT = 16'he4aa;
    SB_LUT4 n12359_bdd_4_lut (.I0(n12359), .I1(ram_s_5_5), .I2(ram_s_4_5), 
            .I3(port_id[1]), .O(n10469));
    defparam n12359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_10670 (.I0(port_id[1]), .I1(n9966), .I2(n9967), 
            .I3(port_id[2]), .O(n11513));
    defparam port_id_1__bdd_4_lut_10670.LUT_INIT = 16'he4aa;
    SB_LUT4 n11939_bdd_4_lut (.I0(n11939), .I1(ram_s_13_5), .I2(ram_s_12_5), 
            .I3(port_id[1]), .O(n11006));
    defparam n11939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1552_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_114_0), .O(n1800));   // src/ram.vhd(68[19:45])
    defparam i1552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11513_bdd_4_lut (.I0(n11513), .I1(n9955), .I2(n9954), .I3(port_id[2]), 
            .O(n11516));
    defparam n11513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10601 (.I0(port_id[0]), .I1(ram_s_42_2), 
            .I2(ram_s_43_2), .I3(port_id[1]), .O(n11747));
    defparam port_id_0__bdd_4_lut_10601.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11095 (.I0(port_id[0]), .I1(ram_s_2_0), 
            .I2(ram_s_3_0), .I3(port_id[1]), .O(n12353));
    defparam port_id_0__bdd_4_lut_11095.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11668 (.I0(port_id[0]), .I1(ram_s_2_1), 
            .I2(ram_s_3_1), .I3(port_id[1]), .O(n13031));
    defparam port_id_0__bdd_4_lut_11668.LUT_INIT = 16'he4aa;
    SB_LUT4 i2535_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_236_7), .O(n2783));   // src/ram.vhd(68[19:45])
    defparam i2535_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12353_bdd_4_lut (.I0(n12353), .I1(ram_s_1_0), .I2(ram_s_0_0), 
            .I3(port_id[1]), .O(n12356));
    defparam n12353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2534_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_236_6), .O(n2782));   // src/ram.vhd(68[19:45])
    defparam i2534_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2533_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_236_5), .O(n2781));   // src/ram.vhd(68[19:45])
    defparam i2533_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10407 (.I0(port_id[0]), .I1(ram_s_66_0), 
            .I2(ram_s_67_0), .I3(port_id[1]), .O(n11507));
    defparam port_id_0__bdd_4_lut_10407.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10910 (.I0(port_id[0]), .I1(ram_s_34_1), 
            .I2(ram_s_35_1), .I3(port_id[1]), .O(n12125));
    defparam port_id_0__bdd_4_lut_10910.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10770 (.I0(port_id[2]), .I1(n9764), .I2(n11606), 
            .I3(port_id[3]), .O(n11933));
    defparam port_id_2__bdd_4_lut_10770.LUT_INIT = 16'he4aa;
    SB_LUT4 n12125_bdd_4_lut (.I0(n12125), .I1(ram_s_33_1), .I2(ram_s_32_1), 
            .I3(port_id[1]), .O(n12128));
    defparam n12125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11933_bdd_4_lut (.I0(n11933), .I1(n9758), .I2(n9740), .I3(port_id[3]), 
            .O(n11009));
    defparam n11933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11219_bdd_4_lut (.I0(n11219), .I1(ram_s_201_1), .I2(ram_s_200_1), 
            .I3(port_id[1]), .O(n11222));
    defparam n11219_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2532_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_236_4), .O(n2780));   // src/ram.vhd(68[19:45])
    defparam i2532_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13031_bdd_4_lut (.I0(n13031), .I1(ram_s_1_1), .I2(ram_s_0_1), 
            .I3(port_id[1]), .O(n13034));
    defparam n13031_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2531_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_236_3), .O(n2779));   // src/ram.vhd(68[19:45])
    defparam i2531_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11507_bdd_4_lut (.I0(n11507), .I1(ram_s_65_0), .I2(ram_s_64_0), 
            .I3(port_id[1]), .O(n11510));
    defparam n11507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11653 (.I0(port_id[0]), .I1(ram_s_10_2), 
            .I2(ram_s_11_2), .I3(port_id[1]), .O(n13025));
    defparam port_id_0__bdd_4_lut_11653.LUT_INIT = 16'he4aa;
    SB_LUT4 n13025_bdd_4_lut (.I0(n13025), .I1(ram_s_9_2), .I2(ram_s_8_2), 
            .I3(port_id[1]), .O(n10808));
    defparam n13025_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10151 (.I0(port_id[0]), .I1(ram_s_146_7), 
            .I2(ram_s_147_7), .I3(port_id[1]), .O(n11213));
    defparam port_id_0__bdd_4_lut_10151.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10387 (.I0(port_id[0]), .I1(ram_s_38_0), 
            .I2(ram_s_39_0), .I3(port_id[1]), .O(n11501));
    defparam port_id_0__bdd_4_lut_10387.LUT_INIT = 16'he4aa;
    SB_LUT4 i2530_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_236_2), .O(n2778));   // src/ram.vhd(68[19:45])
    defparam i2530_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_1__bdd_4_lut_11149 (.I0(port_id[1]), .I1(n10278), .I2(n10279), 
            .I3(port_id[2]), .O(n12347));
    defparam port_id_1__bdd_4_lut_11149.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10900 (.I0(port_id[0]), .I1(ram_s_178_6), 
            .I2(ram_s_179_6), .I3(port_id[1]), .O(n12119));
    defparam port_id_0__bdd_4_lut_10900.LUT_INIT = 16'he4aa;
    SB_LUT4 i2529_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_236_1), .O(n2777));   // src/ram.vhd(68[19:45])
    defparam i2529_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11747_bdd_4_lut (.I0(n11747), .I1(ram_s_41_2), .I2(ram_s_40_2), 
            .I3(port_id[1]), .O(n11750));
    defparam n11747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12119_bdd_4_lut (.I0(n12119), .I1(ram_s_177_6), .I2(ram_s_176_6), 
            .I3(port_id[1]), .O(n12122));
    defparam n12119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11648 (.I0(port_id[0]), .I1(ram_s_114_2), 
            .I2(ram_s_115_2), .I3(port_id[1]), .O(n13019));
    defparam port_id_0__bdd_4_lut_11648.LUT_INIT = 16'he4aa;
    SB_LUT4 n12347_bdd_4_lut (.I0(n12347), .I1(n10264), .I2(n10263), .I3(port_id[2]), 
            .O(n10882));
    defparam n12347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2528_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_236_0), .O(n2776));   // src/ram.vhd(68[19:45])
    defparam i2528_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13019_bdd_4_lut (.I0(n13019), .I1(ram_s_113_2), .I2(ram_s_112_2), 
            .I3(port_id[1]), .O(n13022));
    defparam n13019_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11213_bdd_4_lut (.I0(n11213), .I1(ram_s_145_7), .I2(ram_s_144_7), 
            .I3(port_id[1]), .O(n11216));
    defparam n11213_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11718 (.I0(port_id[2]), .I1(n12032), .I2(n11978), 
            .I3(port_id[3]), .O(n13013));
    defparam port_id_2__bdd_4_lut_11718.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10970 (.I0(port_id[2]), .I1(n11678), .I2(n9116), 
            .I3(port_id[3]), .O(n12113));
    defparam port_id_2__bdd_4_lut_10970.LUT_INIT = 16'he4aa;
    SB_LUT4 n13013_bdd_4_lut (.I0(n13013), .I1(n12068), .I2(n12110), .I3(port_id[3]), 
            .O(n13016));
    defparam n13013_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10740 (.I0(port_id[2]), .I1(n11186), .I2(n9809), 
            .I3(port_id[3]), .O(n11921));
    defparam port_id_2__bdd_4_lut_10740.LUT_INIT = 16'he4aa;
    SB_LUT4 n11921_bdd_4_lut (.I0(n11921), .I1(n11486), .I2(n11600), .I3(port_id[3]), 
            .O(n11015));
    defparam n11921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11643 (.I0(port_id[0]), .I1(ram_s_74_7), 
            .I2(ram_s_75_7), .I3(port_id[1]), .O(n13007));
    defparam port_id_0__bdd_4_lut_11643.LUT_INIT = 16'he4aa;
    SB_LUT4 n12113_bdd_4_lut (.I0(n12113), .I1(n9038), .I2(n9017), .I3(port_id[3]), 
            .O(n12116));
    defparam n12113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13007_bdd_4_lut (.I0(n13007), .I1(ram_s_73_7), .I2(ram_s_72_7), 
            .I3(port_id[1]), .O(n13010));
    defparam n13007_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11090 (.I0(port_id[0]), .I1(ram_s_130_7), 
            .I2(ram_s_131_7), .I3(port_id[1]), .O(n12341));
    defparam port_id_0__bdd_4_lut_11090.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_1__bdd_4_lut_11663 (.I0(port_id[1]), .I1(n9240), .I2(n9241), 
            .I3(port_id[2]), .O(n13001));
    defparam port_id_1__bdd_4_lut_11663.LUT_INIT = 16'he4aa;
    SB_LUT4 i1257_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_77_1), .O(n1505));   // src/ram.vhd(68[19:45])
    defparam i1257_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12341_bdd_4_lut (.I0(n12341), .I1(ram_s_129_7), .I2(ram_s_128_7), 
            .I3(port_id[1]), .O(n12344));
    defparam n12341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10895 (.I0(port_id[0]), .I1(ram_s_18_0), 
            .I2(ram_s_19_0), .I3(port_id[1]), .O(n12107));
    defparam port_id_0__bdd_4_lut_10895.LUT_INIT = 16'he4aa;
    SB_LUT4 i1320_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_85_0), .O(n1568));   // src/ram.vhd(68[19:45])
    defparam i1320_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2335_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_211_7), .O(n2583));   // src/ram.vhd(68[19:45])
    defparam i2335_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1551_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_113_7), .O(n1799));   // src/ram.vhd(68[19:45])
    defparam i1551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11501_bdd_4_lut (.I0(n11501), .I1(ram_s_37_0), .I2(ram_s_36_0), 
            .I3(port_id[1]), .O(n11504));
    defparam n11501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1550_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_113_6), .O(n1798));   // src/ram.vhd(68[19:45])
    defparam i1550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1549_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_113_5), .O(n1797));   // src/ram.vhd(68[19:45])
    defparam i1549_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2334_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_211_6), .O(n2582));   // src/ram.vhd(68[19:45])
    defparam i2334_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2333_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_211_5), .O(n2581));   // src/ram.vhd(68[19:45])
    defparam i2333_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1548_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_113_4), .O(n1796));   // src/ram.vhd(68[19:45])
    defparam i1548_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10586 (.I0(port_id[0]), .I1(ram_s_142_5), 
            .I2(ram_s_143_5), .I3(port_id[1]), .O(n11735));
    defparam port_id_0__bdd_4_lut_10586.LUT_INIT = 16'he4aa;
    SB_LUT4 i1547_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_113_3), .O(n1795));   // src/ram.vhd(68[19:45])
    defparam i1547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12107_bdd_4_lut (.I0(n12107), .I1(ram_s_17_0), .I2(ram_s_16_0), 
            .I3(port_id[1]), .O(n12110));
    defparam n12107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11735_bdd_4_lut (.I0(n11735), .I1(ram_s_141_5), .I2(ram_s_140_5), 
            .I3(port_id[1]), .O(n11738));
    defparam n11735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1546_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_113_2), .O(n1794));   // src/ram.vhd(68[19:45])
    defparam i1546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1545_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_113_1), .O(n1793));   // src/ram.vhd(68[19:45])
    defparam i1545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13001_bdd_4_lut (.I0(n13001), .I1(n9232), .I2(n9231), .I3(port_id[2]), 
            .O(n13004));
    defparam n13001_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11080 (.I0(port_id[0]), .I1(ram_s_30_5), 
            .I2(ram_s_31_5), .I3(port_id[1]), .O(n12335));
    defparam port_id_0__bdd_4_lut_11080.LUT_INIT = 16'he4aa;
    SB_LUT4 i1544_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_113_0), .O(n1792));   // src/ram.vhd(68[19:45])
    defparam i1544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2527_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_235_7), .O(n2775));   // src/ram.vhd(68[19:45])
    defparam i2527_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10576 (.I0(port_id[0]), .I1(ram_s_62_0), 
            .I2(ram_s_63_0), .I3(port_id[1]), .O(n11729));
    defparam port_id_0__bdd_4_lut_10576.LUT_INIT = 16'he4aa;
    SB_LUT4 i2332_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_211_4), .O(n2580));   // src/ram.vhd(68[19:45])
    defparam i2332_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10461 (.I0(port_id[0]), .I1(ram_s_194_1), 
            .I2(ram_s_195_1), .I3(port_id[1]), .O(n11585));
    defparam port_id_0__bdd_4_lut_10461.LUT_INIT = 16'he4aa;
    SB_LUT4 i2526_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_235_6), .O(n2774));   // src/ram.vhd(68[19:45])
    defparam i2526_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12335_bdd_4_lut (.I0(n12335), .I1(ram_s_29_5), .I2(ram_s_28_5), 
            .I3(port_id[1]), .O(n9752));
    defparam n12335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2331_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_211_3), .O(n2579));   // src/ram.vhd(68[19:45])
    defparam i2331_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_2__bdd_4_lut_10730 (.I0(port_id[2]), .I1(n9044), .I2(n9056), 
            .I3(port_id[3]), .O(n11909));
    defparam port_id_2__bdd_4_lut_10730.LUT_INIT = 16'he4aa;
    SB_LUT4 n11729_bdd_4_lut (.I0(n11729), .I1(ram_s_61_0), .I2(ram_s_60_0), 
            .I3(port_id[1]), .O(n11732));
    defparam n11729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2525_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_235_5), .O(n2773));   // src/ram.vhd(68[19:45])
    defparam i2525_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2330_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_211_2), .O(n2578));   // src/ram.vhd(68[19:45])
    defparam i2330_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11585_bdd_4_lut (.I0(n11585), .I1(ram_s_193_1), .I2(ram_s_192_1), 
            .I3(port_id[1]), .O(n11588));
    defparam n11585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2524_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_235_4), .O(n2772));   // src/ram.vhd(68[19:45])
    defparam i2524_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1256_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_77_0), .O(n1504));   // src/ram.vhd(68[19:45])
    defparam i1256_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_1__bdd_4_lut_11628 (.I0(port_id[1]), .I1(n9207), .I2(n9208), 
            .I3(port_id[2]), .O(n12989));
    defparam port_id_1__bdd_4_lut_11628.LUT_INIT = 16'he4aa;
    SB_LUT4 n12989_bdd_4_lut (.I0(n12989), .I1(n9196), .I2(n9195), .I3(port_id[2]), 
            .O(n12992));
    defparam n12989_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11909_bdd_4_lut (.I0(n11909), .I1(n9023), .I2(n9008), .I3(port_id[3]), 
            .O(n11912));
    defparam n11909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11633 (.I0(port_id[0]), .I1(ram_s_74_4), 
            .I2(ram_s_75_4), .I3(port_id[1]), .O(n12983));
    defparam port_id_0__bdd_4_lut_11633.LUT_INIT = 16'he4aa;
    SB_LUT4 n12983_bdd_4_lut (.I0(n12983), .I1(ram_s_73_4), .I2(ram_s_72_4), 
            .I3(port_id[1]), .O(n9692));
    defparam n12983_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10571 (.I0(port_id[0]), .I1(ram_s_42_7), 
            .I2(ram_s_43_7), .I3(port_id[1]), .O(n11723));
    defparam port_id_0__bdd_4_lut_10571.LUT_INIT = 16'he4aa;
    SB_LUT4 n11723_bdd_4_lut (.I0(n11723), .I1(ram_s_41_7), .I2(ram_s_40_7), 
            .I3(port_id[1]), .O(n11726));
    defparam n11723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11618 (.I0(port_id[1]), .I1(n9264), .I2(n9265), 
            .I3(port_id[2]), .O(n12971));
    defparam port_id_1__bdd_4_lut_11618.LUT_INIT = 16'he4aa;
    SB_LUT4 i2523_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_235_3), .O(n2771));   // src/ram.vhd(68[19:45])
    defparam i2523_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10146 (.I0(port_id[0]), .I1(ram_s_74_2), 
            .I2(ram_s_75_2), .I3(port_id[1]), .O(n11207));
    defparam port_id_0__bdd_4_lut_10146.LUT_INIT = 16'he4aa;
    SB_LUT4 i2522_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_235_2), .O(n2770));   // src/ram.vhd(68[19:45])
    defparam i2522_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11207_bdd_4_lut (.I0(n11207), .I1(ram_s_73_2), .I2(ram_s_72_2), 
            .I3(port_id[1]), .O(n11210));
    defparam n11207_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2521_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_235_1), .O(n2769));   // src/ram.vhd(68[19:45])
    defparam i2521_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2520_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_235_0), .O(n2768));   // src/ram.vhd(68[19:45])
    defparam i2520_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_2__bdd_4_lut_10170 (.I0(port_id[2]), .I1(n9794), .I2(n9818), 
            .I3(port_id[3]), .O(n11201));
    defparam port_id_2__bdd_4_lut_10170.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10451 (.I0(port_id[0]), .I1(ram_s_86_7), 
            .I2(ram_s_87_7), .I3(port_id[1]), .O(n11579));
    defparam port_id_0__bdd_4_lut_10451.LUT_INIT = 16'he4aa;
    SB_LUT4 n11201_bdd_4_lut (.I0(n11201), .I1(n9746), .I2(n9725), .I3(port_id[3]), 
            .O(n11204));
    defparam n11201_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2519_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_234_7), .O(n2767));   // src/ram.vhd(68[19:45])
    defparam i2519_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2303_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_207_7), .O(n2551));   // src/ram.vhd(68[19:45])
    defparam i2303_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2518_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_234_6), .O(n2766));   // src/ram.vhd(68[19:45])
    defparam i2518_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2517_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_234_5), .O(n2765));   // src/ram.vhd(68[19:45])
    defparam i2517_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12971_bdd_4_lut (.I0(n12971), .I1(n9253), .I2(n9252), .I3(port_id[2]), 
            .O(n12974));
    defparam n12971_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2329_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_211_1), .O(n2577));   // src/ram.vhd(68[19:45])
    defparam i2329_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2516_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_234_4), .O(n2764));   // src/ram.vhd(68[19:45])
    defparam i2516_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11613 (.I0(port_id[0]), .I1(ram_s_186_3), 
            .I2(ram_s_187_3), .I3(port_id[1]), .O(n12965));
    defparam port_id_0__bdd_4_lut_11613.LUT_INIT = 16'he4aa;
    SB_LUT4 n12965_bdd_4_lut (.I0(n12965), .I1(ram_s_185_3), .I2(ram_s_184_3), 
            .I3(port_id[1]), .O(n12968));
    defparam n12965_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11603 (.I0(port_id[1]), .I1(n9171), .I2(n9172), 
            .I3(port_id[2]), .O(n12959));
    defparam port_id_1__bdd_4_lut_11603.LUT_INIT = 16'he4aa;
    SB_LUT4 n12959_bdd_4_lut (.I0(n12959), .I1(n9163), .I2(n9162), .I3(port_id[2]), 
            .O(n12962));
    defparam n12959_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1248_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_76_0), .O(n1496));   // src/ram.vhd(68[19:45])
    defparam i1248_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2302_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_207_6), .O(n2550));   // src/ram.vhd(68[19:45])
    defparam i2302_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10885 (.I0(port_id[0]), .I1(ram_s_206_7), 
            .I2(ram_s_207_7), .I3(port_id[1]), .O(n12095));
    defparam port_id_0__bdd_4_lut_10885.LUT_INIT = 16'he4aa;
    SB_LUT4 n11579_bdd_4_lut (.I0(n11579), .I1(ram_s_85_7), .I2(ram_s_84_7), 
            .I3(port_id[1]), .O(n11582));
    defparam n11579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11638 (.I0(port_id[2]), .I1(n10634), .I2(n10649), 
            .I3(port_id[3]), .O(n12953));
    defparam port_id_2__bdd_4_lut_11638.LUT_INIT = 16'he4aa;
    SB_LUT4 n12953_bdd_4_lut (.I0(n12953), .I1(n10625), .I2(n10622), .I3(port_id[3]), 
            .O(n10811));
    defparam n12953_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10566 (.I0(port_id[0]), .I1(ram_s_214_7), 
            .I2(ram_s_215_7), .I3(port_id[1]), .O(n11717));
    defparam port_id_0__bdd_4_lut_10566.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11075 (.I0(port_id[0]), .I1(ram_s_190_2), 
            .I2(ram_s_191_2), .I3(port_id[1]), .O(n12329));
    defparam port_id_0__bdd_4_lut_11075.LUT_INIT = 16'he4aa;
    SB_LUT4 n12095_bdd_4_lut (.I0(n12095), .I1(ram_s_205_7), .I2(ram_s_204_7), 
            .I3(port_id[1]), .O(n10499));
    defparam n12095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11717_bdd_4_lut (.I0(n11717), .I1(ram_s_213_7), .I2(ram_s_212_7), 
            .I3(port_id[1]), .O(n10532));
    defparam n11717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2515_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_234_3), .O(n2763));   // src/ram.vhd(68[19:45])
    defparam i2515_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10446 (.I0(port_id[0]), .I1(ram_s_42_1), 
            .I2(ram_s_43_1), .I3(port_id[1]), .O(n11573));
    defparam port_id_0__bdd_4_lut_10446.LUT_INIT = 16'he4aa;
    SB_LUT4 i2514_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_234_2), .O(n2762));   // src/ram.vhd(68[19:45])
    defparam i2514_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2328_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_211_0), .O(n2576));   // src/ram.vhd(68[19:45])
    defparam i2328_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i174_2_lut_3_lut (.I0(n45), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n174));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i174_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i2513_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_234_1), .O(n2761));   // src/ram.vhd(68[19:45])
    defparam i2513_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2512_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_234_0), .O(n2760));   // src/ram.vhd(68[19:45])
    defparam i2512_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1543_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_112_7), .O(n1791));   // src/ram.vhd(68[19:45])
    defparam i1543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1542_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_112_6), .O(n1790));   // src/ram.vhd(68[19:45])
    defparam i1542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1541_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_112_5), .O(n1789));   // src/ram.vhd(68[19:45])
    defparam i1541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1540_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_112_4), .O(n1788));   // src/ram.vhd(68[19:45])
    defparam i1540_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11573_bdd_4_lut (.I0(n11573), .I1(ram_s_41_1), .I2(ram_s_40_1), 
            .I3(port_id[1]), .O(n11576));
    defparam n11573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1539_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_112_3), .O(n1787));   // src/ram.vhd(68[19:45])
    defparam i1539_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1538_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_112_2), .O(n1786));   // src/ram.vhd(68[19:45])
    defparam i1538_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1537_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_112_1), .O(n1785));   // src/ram.vhd(68[19:45])
    defparam i1537_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1536_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_112_0), .O(n1784));   // src/ram.vhd(68[19:45])
    defparam i1536_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2511_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_233_7), .O(n2759));   // src/ram.vhd(68[19:45])
    defparam i2511_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2510_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_233_6), .O(n2758));   // src/ram.vhd(68[19:45])
    defparam i2510_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2509_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_233_5), .O(n2757));   // src/ram.vhd(68[19:45])
    defparam i2509_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2508_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_233_4), .O(n2756));   // src/ram.vhd(68[19:45])
    defparam i2508_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10561 (.I0(port_id[0]), .I1(ram_s_6_7), 
            .I2(ram_s_7_7), .I3(port_id[1]), .O(n11711));
    defparam port_id_0__bdd_4_lut_10561.LUT_INIT = 16'he4aa;
    SB_LUT4 i2507_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_233_3), .O(n2755));   // src/ram.vhd(68[19:45])
    defparam i2507_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11598 (.I0(port_id[0]), .I1(ram_s_134_0), 
            .I2(ram_s_135_0), .I3(port_id[1]), .O(n12947));
    defparam port_id_0__bdd_4_lut_11598.LUT_INIT = 16'he4aa;
    SB_LUT4 n11711_bdd_4_lut (.I0(n11711), .I1(ram_s_5_7), .I2(ram_s_4_7), 
            .I3(port_id[1]), .O(n11714));
    defparam n11711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12947_bdd_4_lut (.I0(n12947), .I1(ram_s_133_0), .I2(ram_s_132_0), 
            .I3(port_id[1]), .O(n9065));
    defparam n12947_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12329_bdd_4_lut (.I0(n12329), .I1(ram_s_189_2), .I2(ram_s_188_2), 
            .I3(port_id[1]), .O(n12332));
    defparam n12329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10875 (.I0(port_id[0]), .I1(ram_s_34_2), 
            .I2(ram_s_35_2), .I3(port_id[1]), .O(n12089));
    defparam port_id_0__bdd_4_lut_10875.LUT_INIT = 16'he4aa;
    SB_LUT4 i2506_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_233_2), .O(n2754));   // src/ram.vhd(68[19:45])
    defparam i2506_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i173_2_lut_3_lut (.I0(n45), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n173));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i173_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2505_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_233_1), .O(n2753));   // src/ram.vhd(68[19:45])
    defparam i2505_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1319_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_84_7), .O(n1567));   // src/ram.vhd(68[19:45])
    defparam i1319_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1318_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_84_6), .O(n1566));   // src/ram.vhd(68[19:45])
    defparam i1318_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1317_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_84_5), .O(n1565));   // src/ram.vhd(68[19:45])
    defparam i1317_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1316_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_84_4), .O(n1564));   // src/ram.vhd(68[19:45])
    defparam i1316_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1315_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_84_3), .O(n1563));   // src/ram.vhd(68[19:45])
    defparam i1315_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1314_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_84_2), .O(n1562));   // src/ram.vhd(68[19:45])
    defparam i1314_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1313_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_84_1), .O(n1561));   // src/ram.vhd(68[19:45])
    defparam i1313_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1312_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_84_0), .O(n1560));   // src/ram.vhd(68[19:45])
    defparam i1312_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_1__bdd_4_lut_11593 (.I0(port_id[1]), .I1(n9855), .I2(n9856), 
            .I3(port_id[2]), .O(n12941));
    defparam port_id_1__bdd_4_lut_11593.LUT_INIT = 16'he4aa;
    SB_LUT4 i2504_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_233_0), .O(n2752));   // src/ram.vhd(68[19:45])
    defparam i2504_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12941_bdd_4_lut (.I0(n12941), .I1(n9814), .I2(n9813), .I3(port_id[2]), 
            .O(n10813));
    defparam n12941_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1535_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_111_7), .O(n1783));   // src/ram.vhd(68[19:45])
    defparam i1535_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10556 (.I0(port_id[0]), .I1(ram_s_58_5), 
            .I2(ram_s_59_5), .I3(port_id[1]), .O(n11705));
    defparam port_id_0__bdd_4_lut_10556.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_1__bdd_4_lut_11578 (.I0(port_id[1]), .I1(n9141), .I2(n9142), 
            .I3(port_id[2]), .O(n12935));
    defparam port_id_1__bdd_4_lut_11578.LUT_INIT = 16'he4aa;
    SB_LUT4 i2327_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_210_7), .O(n2575));   // src/ram.vhd(68[19:45])
    defparam i2327_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1534_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_111_6), .O(n1782));   // src/ram.vhd(68[19:45])
    defparam i1534_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12935_bdd_4_lut (.I0(n12935), .I1(n9127), .I2(n9126), .I3(port_id[2]), 
            .O(n12938));
    defparam n12935_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11583 (.I0(port_id[0]), .I1(ram_s_182_2), 
            .I2(ram_s_183_2), .I3(port_id[1]), .O(n12929));
    defparam port_id_0__bdd_4_lut_11583.LUT_INIT = 16'he4aa;
    SB_LUT4 n12929_bdd_4_lut (.I0(n12929), .I1(ram_s_181_2), .I2(ram_s_180_2), 
            .I3(port_id[1]), .O(n12932));
    defparam n12929_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1533_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_111_5), .O(n1781));   // src/ram.vhd(68[19:45])
    defparam i1533_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1532_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_111_4), .O(n1780));   // src/ram.vhd(68[19:45])
    defparam i1532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1531_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_111_3), .O(n1779));   // src/ram.vhd(68[19:45])
    defparam i1531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1530_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_111_2), .O(n1778));   // src/ram.vhd(68[19:45])
    defparam i1530_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1529_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_111_1), .O(n1777));   // src/ram.vhd(68[19:45])
    defparam i1529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1528_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_111_0), .O(n1776));   // src/ram.vhd(68[19:45])
    defparam i1528_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10141 (.I0(port_id[0]), .I1(ram_s_50_0), 
            .I2(ram_s_51_0), .I3(port_id[1]), .O(n11195));
    defparam port_id_0__bdd_4_lut_10141.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10516 (.I0(port_id[2]), .I1(n10541), .I2(n11252), 
            .I3(port_id[3]), .O(n11567));
    defparam port_id_2__bdd_4_lut_10516.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11568 (.I0(port_id[0]), .I1(ram_s_58_0), 
            .I2(ram_s_59_0), .I3(port_id[1]), .O(n12917));
    defparam port_id_0__bdd_4_lut_11568.LUT_INIT = 16'he4aa;
    SB_LUT4 n12917_bdd_4_lut (.I0(n12917), .I1(ram_s_57_0), .I2(ram_s_56_0), 
            .I3(port_id[1]), .O(n8906));
    defparam n12917_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11558 (.I0(port_id[0]), .I1(ram_s_94_5), 
            .I2(ram_s_95_5), .I3(port_id[1]), .O(n12911));
    defparam port_id_0__bdd_4_lut_11558.LUT_INIT = 16'he4aa;
    SB_LUT4 n12911_bdd_4_lut (.I0(n12911), .I1(ram_s_93_5), .I2(ram_s_92_5), 
            .I3(port_id[1]), .O(n12914));
    defparam n12911_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11588 (.I0(port_id[2]), .I1(n10808), .I2(n12698), 
            .I3(port_id[3]), .O(n12905));
    defparam port_id_2__bdd_4_lut_11588.LUT_INIT = 16'he4aa;
    SB_LUT4 n12905_bdd_4_lut (.I0(n12905), .I1(n10796), .I2(n10772), .I3(port_id[3]), 
            .O(n12908));
    defparam n12905_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11553 (.I0(port_id[0]), .I1(ram_s_138_0), 
            .I2(ram_s_139_0), .I3(port_id[1]), .O(n12899));
    defparam port_id_0__bdd_4_lut_11553.LUT_INIT = 16'he4aa;
    SB_LUT4 n12899_bdd_4_lut (.I0(n12899), .I1(ram_s_137_0), .I2(ram_s_136_0), 
            .I3(port_id[1]), .O(n9068));
    defparam n12899_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11573 (.I0(port_id[1]), .I1(n9135), .I2(n9136), 
            .I3(port_id[2]), .O(n12893));
    defparam port_id_1__bdd_4_lut_11573.LUT_INIT = 16'he4aa;
    SB_LUT4 i2326_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_210_6), .O(n2574));   // src/ram.vhd(68[19:45])
    defparam i2326_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2503_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_232_7), .O(n2751));   // src/ram.vhd(68[19:45])
    defparam i2503_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2502_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_232_6), .O(n2750));   // src/ram.vhd(68[19:45])
    defparam i2502_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11567_bdd_4_lut (.I0(n11567), .I1(n10532), .I2(n10517), .I3(port_id[3]), 
            .O(n11570));
    defparam n11567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12893_bdd_4_lut (.I0(n12893), .I1(n9061), .I2(n9060), .I3(port_id[2]), 
            .O(n10816));
    defparam n12893_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11543 (.I0(port_id[0]), .I1(ram_s_190_5), 
            .I2(ram_s_191_5), .I3(port_id[1]), .O(n12887));
    defparam port_id_0__bdd_4_lut_11543.LUT_INIT = 16'he4aa;
    SB_LUT4 n12887_bdd_4_lut (.I0(n12887), .I1(ram_s_189_5), .I2(ram_s_188_5), 
            .I3(port_id[1]), .O(n9701));
    defparam n12887_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11548 (.I0(port_id[2]), .I1(n11456), .I2(n11288), 
            .I3(port_id[3]), .O(n12881));
    defparam port_id_2__bdd_4_lut_11548.LUT_INIT = 16'he4aa;
    SB_LUT4 n12881_bdd_4_lut (.I0(n12881), .I1(n11504), .I2(n11774), .I3(port_id[3]), 
            .O(n12884));
    defparam n12881_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11533 (.I0(port_id[0]), .I1(ram_s_250_4), 
            .I2(ram_s_251_4), .I3(port_id[1]), .O(n12875));
    defparam port_id_0__bdd_4_lut_11533.LUT_INIT = 16'he4aa;
    SB_LUT4 i2501_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_232_5), .O(n2749));   // src/ram.vhd(68[19:45])
    defparam i2501_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2500_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_232_4), .O(n2748));   // src/ram.vhd(68[19:45])
    defparam i2500_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12875_bdd_4_lut (.I0(n12875), .I1(ram_s_249_4), .I2(ram_s_248_4), 
            .I3(port_id[1]), .O(n12878));
    defparam n12875_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11528 (.I0(port_id[2]), .I1(n8906), .I2(n11732), 
            .I3(port_id[3]), .O(n12869));
    defparam port_id_2__bdd_4_lut_11528.LUT_INIT = 16'he4aa;
    SB_LUT4 n11705_bdd_4_lut (.I0(n11705), .I1(ram_s_57_5), .I2(ram_s_56_5), 
            .I3(port_id[1]), .O(n11708));
    defparam n11705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12089_bdd_4_lut (.I0(n12089), .I1(ram_s_33_2), .I2(ram_s_32_2), 
            .I3(port_id[1]), .O(n12092));
    defparam n12089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10720 (.I0(port_id[2]), .I1(n9872), .I2(n9881), 
            .I3(port_id[3]), .O(n11891));
    defparam port_id_2__bdd_4_lut_10720.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10441 (.I0(port_id[0]), .I1(ram_s_142_7), 
            .I2(ram_s_143_7), .I3(port_id[1]), .O(n11561));
    defparam port_id_0__bdd_4_lut_10441.LUT_INIT = 16'he4aa;
    SB_LUT4 i2325_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_210_5), .O(n2573));   // src/ram.vhd(68[19:45])
    defparam i2325_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11891_bdd_4_lut (.I0(n11891), .I1(n9863), .I2(n9854), .I3(port_id[3]), 
            .O(n11033));
    defparam n11891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12869_bdd_4_lut (.I0(n12869), .I1(n11966), .I2(n11198), .I3(port_id[3]), 
            .O(n12872));
    defparam n12869_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11561_bdd_4_lut (.I0(n11561), .I1(ram_s_141_7), .I2(ram_s_140_7), 
            .I3(port_id[1]), .O(n11564));
    defparam n11561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11070 (.I0(port_id[0]), .I1(ram_s_110_3), 
            .I2(ram_s_111_3), .I3(port_id[1]), .O(n12323));
    defparam port_id_0__bdd_4_lut_11070.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10551 (.I0(port_id[0]), .I1(ram_s_94_6), 
            .I2(ram_s_95_6), .I3(port_id[1]), .O(n11699));
    defparam port_id_0__bdd_4_lut_10551.LUT_INIT = 16'he4aa;
    SB_LUT4 n12323_bdd_4_lut (.I0(n12323), .I1(ram_s_109_3), .I2(ram_s_108_3), 
            .I3(port_id[1]), .O(n9395));
    defparam n12323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11699_bdd_4_lut (.I0(n11699), .I1(ram_s_93_6), .I2(ram_s_92_6), 
            .I3(port_id[1]), .O(n11702));
    defparam n11699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11523 (.I0(port_id[0]), .I1(ram_s_82_5), 
            .I2(ram_s_83_5), .I3(port_id[1]), .O(n12863));
    defparam port_id_0__bdd_4_lut_11523.LUT_INIT = 16'he4aa;
    SB_LUT4 n12863_bdd_4_lut (.I0(n12863), .I1(ram_s_81_5), .I2(ram_s_80_5), 
            .I3(port_id[1]), .O(n12866));
    defparam n12863_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2499_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_232_3), .O(n2747));   // src/ram.vhd(68[19:45])
    defparam i2499_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11065 (.I0(port_id[0]), .I1(ram_s_158_1), 
            .I2(ram_s_159_1), .I3(port_id[1]), .O(n12317));
    defparam port_id_0__bdd_4_lut_11065.LUT_INIT = 16'he4aa;
    SB_LUT4 n12317_bdd_4_lut (.I0(n12317), .I1(ram_s_157_1), .I2(ram_s_156_1), 
            .I3(port_id[1]), .O(n12320));
    defparam n12317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10546 (.I0(port_id[0]), .I1(ram_s_190_1), 
            .I2(ram_s_191_1), .I3(port_id[1]), .O(n11693));
    defparam port_id_0__bdd_4_lut_10546.LUT_INIT = 16'he4aa;
    SB_LUT4 n11195_bdd_4_lut (.I0(n11195), .I1(ram_s_49_0), .I2(ram_s_48_0), 
            .I3(port_id[1]), .O(n11198));
    defparam n11195_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i248_249 (.Q(ram_s_9_6), .C(CLK_3P3_MHZ_c), .D(n897));   // src/ram.vhd(56[12:17])
    SB_LUT4 port_id_0__bdd_4_lut_11513 (.I0(port_id[0]), .I1(ram_s_138_1), 
            .I2(ram_s_139_1), .I3(port_id[1]), .O(n12857));
    defparam port_id_0__bdd_4_lut_11513.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10705 (.I0(port_id[2]), .I1(n9662), .I2(n9671), 
            .I3(port_id[3]), .O(n11885));
    defparam port_id_2__bdd_4_lut_10705.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_1__bdd_4_lut_10180 (.I0(port_id[1]), .I1(n9999), .I2(n10000), 
            .I3(port_id[2]), .O(n11189));
    defparam port_id_1__bdd_4_lut_10180.LUT_INIT = 16'he4aa;
    SB_LUT4 n11885_bdd_4_lut (.I0(n11885), .I1(n9644), .I2(n9635), .I3(port_id[3]), 
            .O(n11888));
    defparam n11885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12857_bdd_4_lut (.I0(n12857), .I1(ram_s_137_1), .I2(ram_s_136_1), 
            .I3(port_id[1]), .O(n12860));
    defparam n12857_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i254_255 (.Q(ram_s_10_0), .C(CLK_3P3_MHZ_c), .D(n896));   // src/ram.vhd(56[12:17])
    SB_DFF i263_264 (.Q(ram_s_10_3), .C(CLK_3P3_MHZ_c), .D(n895));   // src/ram.vhd(56[12:17])
    SB_LUT4 port_id_0__bdd_4_lut_11508 (.I0(port_id[0]), .I1(ram_s_38_7), 
            .I2(ram_s_39_7), .I3(port_id[1]), .O(n12851));
    defparam port_id_0__bdd_4_lut_11508.LUT_INIT = 16'he4aa;
    SB_DFF i257_258 (.Q(ram_s_10_1), .C(CLK_3P3_MHZ_c), .D(n894));   // src/ram.vhd(56[12:17])
    SB_LUT4 n12851_bdd_4_lut (.I0(n12851), .I1(ram_s_37_7), .I2(ram_s_36_7), 
            .I3(port_id[1]), .O(n12854));
    defparam n12851_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11189_bdd_4_lut (.I0(n11189), .I1(n9991), .I2(n9990), .I3(port_id[2]), 
            .O(n11192));
    defparam n11189_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i362_363 (.Q(ram_s_14_4), .C(CLK_3P3_MHZ_c), .D(n893));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2498_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_232_2), .O(n2746));   // src/ram.vhd(68[19:45])
    defparam i2498_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11503 (.I0(port_id[0]), .I1(ram_s_250_6), 
            .I2(ram_s_251_6), .I3(port_id[1]), .O(n12845));
    defparam port_id_0__bdd_4_lut_11503.LUT_INIT = 16'he4aa;
    SB_DFF i527_528 (.Q(ram_s_21_3), .C(CLK_3P3_MHZ_c), .D(n892));   // src/ram.vhd(56[12:17])
    SB_LUT4 n12845_bdd_4_lut (.I0(n12845), .I1(ram_s_249_6), .I2(ram_s_248_6), 
            .I3(port_id[1]), .O(n12848));
    defparam n12845_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i422_423 (.Q(ram_s_17_0), .C(CLK_3P3_MHZ_c), .D(n891));   // src/ram.vhd(56[12:17])
    SB_DFF i425_426 (.Q(ram_s_17_1), .C(CLK_3P3_MHZ_c), .D(n890));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2497_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_232_1), .O(n2745));   // src/ram.vhd(68[19:45])
    defparam i2497_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11498 (.I0(port_id[0]), .I1(ram_s_78_4), 
            .I2(ram_s_79_4), .I3(port_id[1]), .O(n12839));
    defparam port_id_0__bdd_4_lut_11498.LUT_INIT = 16'he4aa;
    SB_DFF i428_429 (.Q(ram_s_17_2), .C(CLK_3P3_MHZ_c), .D(n889));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2496_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_232_0), .O(n2744));   // src/ram.vhd(68[19:45])
    defparam i2496_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12839_bdd_4_lut (.I0(n12839), .I1(ram_s_77_4), .I2(ram_s_76_4), 
            .I3(port_id[1]), .O(n9707));
    defparam n12839_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2324_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_210_4), .O(n2572));   // src/ram.vhd(68[19:45])
    defparam i2324_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i431_432 (.Q(ram_s_17_3), .C(CLK_3P3_MHZ_c), .D(n888));   // src/ram.vhd(56[12:17])
    SB_LUT4 port_id_0__bdd_4_lut_11493 (.I0(port_id[0]), .I1(ram_s_190_7), 
            .I2(ram_s_191_7), .I3(port_id[1]), .O(n12833));
    defparam port_id_0__bdd_4_lut_11493.LUT_INIT = 16'he4aa;
    SB_LUT4 n12833_bdd_4_lut (.I0(n12833), .I1(ram_s_189_7), .I2(ram_s_188_7), 
            .I3(port_id[1]), .O(n10427));
    defparam n12833_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10382 (.I0(port_id[0]), .I1(ram_s_118_4), 
            .I2(ram_s_119_4), .I3(port_id[1]), .O(n11483));
    defparam port_id_0__bdd_4_lut_10382.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10132 (.I0(port_id[0]), .I1(ram_s_122_4), 
            .I2(ram_s_123_4), .I3(port_id[1]), .O(n11183));
    defparam port_id_0__bdd_4_lut_10132.LUT_INIT = 16'he4aa;
    SB_LUT4 n11483_bdd_4_lut (.I0(n11483), .I1(ram_s_117_4), .I2(ram_s_116_4), 
            .I3(port_id[1]), .O(n11486));
    defparam n11483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10367 (.I0(port_id[0]), .I1(ram_s_46_2), 
            .I2(ram_s_47_2), .I3(port_id[1]), .O(n11477));
    defparam port_id_0__bdd_4_lut_10367.LUT_INIT = 16'he4aa;
    SB_LUT4 i1527_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_110_7), .O(n1775));   // src/ram.vhd(68[19:45])
    defparam i1527_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i434_435 (.Q(ram_s_17_4), .C(CLK_3P3_MHZ_c), .D(n887));   // src/ram.vhd(56[12:17])
    SB_DFF i266_267 (.Q(ram_s_10_4), .C(CLK_3P3_MHZ_c), .D(n886));   // src/ram.vhd(56[12:17])
    SB_DFF i437_438 (.Q(ram_s_17_5), .C(CLK_3P3_MHZ_c), .D(n885));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1526_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_110_6), .O(n1774));   // src/ram.vhd(68[19:45])
    defparam i1526_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11477_bdd_4_lut (.I0(n11477), .I1(ram_s_45_2), .I2(ram_s_44_2), 
            .I3(port_id[1]), .O(n11480));
    defparam n11477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1525_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_110_5), .O(n1773));   // src/ram.vhd(68[19:45])
    defparam i1525_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1524_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_110_4), .O(n1772));   // src/ram.vhd(68[19:45])
    defparam i1524_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1523_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_110_3), .O(n1771));   // src/ram.vhd(68[19:45])
    defparam i1523_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1522_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_110_2), .O(n1770));   // src/ram.vhd(68[19:45])
    defparam i1522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1521_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_110_1), .O(n1769));   // src/ram.vhd(68[19:45])
    defparam i1521_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1520_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_110_0), .O(n1768));   // src/ram.vhd(68[19:45])
    defparam i1520_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2495_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_231_7), .O(n2743));   // src/ram.vhd(68[19:45])
    defparam i2495_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2323_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_210_3), .O(n2571));   // src/ram.vhd(68[19:45])
    defparam i2323_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11488 (.I0(port_id[0]), .I1(ram_s_134_5), 
            .I2(ram_s_135_5), .I3(port_id[1]), .O(n12827));
    defparam port_id_0__bdd_4_lut_11488.LUT_INIT = 16'he4aa;
    SB_LUT4 n11183_bdd_4_lut (.I0(n11183), .I1(ram_s_121_4), .I2(ram_s_120_4), 
            .I3(port_id[1]), .O(n11186));
    defparam n11183_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12827_bdd_4_lut (.I0(n12827), .I1(ram_s_133_5), .I2(ram_s_132_5), 
            .I3(port_id[1]), .O(n12830));
    defparam n12827_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2494_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_231_6), .O(n2742));   // src/ram.vhd(68[19:45])
    defparam i2494_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2493_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_231_5), .O(n2741));   // src/ram.vhd(68[19:45])
    defparam i2493_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2492_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_231_4), .O(n2740));   // src/ram.vhd(68[19:45])
    defparam i2492_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i6155_6156 (.Q(ram_s_255_7), .C(CLK_3P3_MHZ_c), .D(n2935));   // src/ram.vhd(56[12:17])
    SB_DFF i6152_6153 (.Q(ram_s_255_6), .C(CLK_3P3_MHZ_c), .D(n2934));   // src/ram.vhd(56[12:17])
    SB_DFF i6149_6150 (.Q(ram_s_255_5), .C(CLK_3P3_MHZ_c), .D(n2933));   // src/ram.vhd(56[12:17])
    SB_DFF i6146_6147 (.Q(ram_s_255_4), .C(CLK_3P3_MHZ_c), .D(n2932));   // src/ram.vhd(56[12:17])
    SB_DFF i6143_6144 (.Q(ram_s_255_3), .C(CLK_3P3_MHZ_c), .D(n2931));   // src/ram.vhd(56[12:17])
    SB_DFF i6140_6141 (.Q(ram_s_255_2), .C(CLK_3P3_MHZ_c), .D(n2930));   // src/ram.vhd(56[12:17])
    SB_DFF i6137_6138 (.Q(ram_s_255_1), .C(CLK_3P3_MHZ_c), .D(n2929));   // src/ram.vhd(56[12:17])
    SB_DFF i6134_6135 (.Q(ram_s_255_0), .C(CLK_3P3_MHZ_c), .D(n2928));   // src/ram.vhd(56[12:17])
    SB_DFF i6131_6132 (.Q(ram_s_254_7), .C(CLK_3P3_MHZ_c), .D(n2927));   // src/ram.vhd(56[12:17])
    SB_DFF i6128_6129 (.Q(ram_s_254_6), .C(CLK_3P3_MHZ_c), .D(n2926));   // src/ram.vhd(56[12:17])
    SB_DFF i6125_6126 (.Q(ram_s_254_5), .C(CLK_3P3_MHZ_c), .D(n2925));   // src/ram.vhd(56[12:17])
    SB_DFF i6122_6123 (.Q(ram_s_254_4), .C(CLK_3P3_MHZ_c), .D(n2924));   // src/ram.vhd(56[12:17])
    SB_DFF i6119_6120 (.Q(ram_s_254_3), .C(CLK_3P3_MHZ_c), .D(n2923));   // src/ram.vhd(56[12:17])
    SB_DFF i6116_6117 (.Q(ram_s_254_2), .C(CLK_3P3_MHZ_c), .D(n2922));   // src/ram.vhd(56[12:17])
    SB_DFF i6113_6114 (.Q(ram_s_254_1), .C(CLK_3P3_MHZ_c), .D(n2921));   // src/ram.vhd(56[12:17])
    SB_DFF i6110_6111 (.Q(ram_s_254_0), .C(CLK_3P3_MHZ_c), .D(n2920));   // src/ram.vhd(56[12:17])
    SB_DFF i6107_6108 (.Q(ram_s_253_7), .C(CLK_3P3_MHZ_c), .D(n2919));   // src/ram.vhd(56[12:17])
    SB_DFF i6104_6105 (.Q(ram_s_253_6), .C(CLK_3P3_MHZ_c), .D(n2918));   // src/ram.vhd(56[12:17])
    SB_DFF i6101_6102 (.Q(ram_s_253_5), .C(CLK_3P3_MHZ_c), .D(n2917));   // src/ram.vhd(56[12:17])
    SB_DFF i6098_6099 (.Q(ram_s_253_4), .C(CLK_3P3_MHZ_c), .D(n2916));   // src/ram.vhd(56[12:17])
    SB_DFF i6095_6096 (.Q(ram_s_253_3), .C(CLK_3P3_MHZ_c), .D(n2915));   // src/ram.vhd(56[12:17])
    SB_DFF i6092_6093 (.Q(ram_s_253_2), .C(CLK_3P3_MHZ_c), .D(n2914));   // src/ram.vhd(56[12:17])
    SB_DFF i6089_6090 (.Q(ram_s_253_1), .C(CLK_3P3_MHZ_c), .D(n2913));   // src/ram.vhd(56[12:17])
    SB_DFF i6086_6087 (.Q(ram_s_253_0), .C(CLK_3P3_MHZ_c), .D(n2912));   // src/ram.vhd(56[12:17])
    SB_DFF i6083_6084 (.Q(ram_s_252_7), .C(CLK_3P3_MHZ_c), .D(n2911));   // src/ram.vhd(56[12:17])
    SB_DFF i6080_6081 (.Q(ram_s_252_6), .C(CLK_3P3_MHZ_c), .D(n2910));   // src/ram.vhd(56[12:17])
    SB_DFF i6077_6078 (.Q(ram_s_252_5), .C(CLK_3P3_MHZ_c), .D(n2909));   // src/ram.vhd(56[12:17])
    SB_DFF i6074_6075 (.Q(ram_s_252_4), .C(CLK_3P3_MHZ_c), .D(n2908));   // src/ram.vhd(56[12:17])
    SB_DFF i6071_6072 (.Q(ram_s_252_3), .C(CLK_3P3_MHZ_c), .D(n2907));   // src/ram.vhd(56[12:17])
    SB_DFF i6068_6069 (.Q(ram_s_252_2), .C(CLK_3P3_MHZ_c), .D(n2906));   // src/ram.vhd(56[12:17])
    SB_DFF i6065_6066 (.Q(ram_s_252_1), .C(CLK_3P3_MHZ_c), .D(n2905));   // src/ram.vhd(56[12:17])
    SB_DFF i6062_6063 (.Q(ram_s_252_0), .C(CLK_3P3_MHZ_c), .D(n2904));   // src/ram.vhd(56[12:17])
    SB_DFF i6059_6060 (.Q(ram_s_251_7), .C(CLK_3P3_MHZ_c), .D(n2903));   // src/ram.vhd(56[12:17])
    SB_DFF i6056_6057 (.Q(ram_s_251_6), .C(CLK_3P3_MHZ_c), .D(n2902));   // src/ram.vhd(56[12:17])
    SB_DFF i6053_6054 (.Q(ram_s_251_5), .C(CLK_3P3_MHZ_c), .D(n2901));   // src/ram.vhd(56[12:17])
    SB_DFF i6050_6051 (.Q(ram_s_251_4), .C(CLK_3P3_MHZ_c), .D(n2900));   // src/ram.vhd(56[12:17])
    SB_DFF i6047_6048 (.Q(ram_s_251_3), .C(CLK_3P3_MHZ_c), .D(n2899));   // src/ram.vhd(56[12:17])
    SB_DFF i6044_6045 (.Q(ram_s_251_2), .C(CLK_3P3_MHZ_c), .D(n2898));   // src/ram.vhd(56[12:17])
    SB_DFF i6041_6042 (.Q(ram_s_251_1), .C(CLK_3P3_MHZ_c), .D(n2897));   // src/ram.vhd(56[12:17])
    SB_DFF i6038_6039 (.Q(ram_s_251_0), .C(CLK_3P3_MHZ_c), .D(n2896));   // src/ram.vhd(56[12:17])
    SB_DFF i6035_6036 (.Q(ram_s_250_7), .C(CLK_3P3_MHZ_c), .D(n2895));   // src/ram.vhd(56[12:17])
    SB_DFF i6032_6033 (.Q(ram_s_250_6), .C(CLK_3P3_MHZ_c), .D(n2894));   // src/ram.vhd(56[12:17])
    SB_DFF i6029_6030 (.Q(ram_s_250_5), .C(CLK_3P3_MHZ_c), .D(n2893));   // src/ram.vhd(56[12:17])
    SB_DFF i6026_6027 (.Q(ram_s_250_4), .C(CLK_3P3_MHZ_c), .D(n2892));   // src/ram.vhd(56[12:17])
    SB_DFF i6023_6024 (.Q(ram_s_250_3), .C(CLK_3P3_MHZ_c), .D(n2891));   // src/ram.vhd(56[12:17])
    SB_DFF i6020_6021 (.Q(ram_s_250_2), .C(CLK_3P3_MHZ_c), .D(n2890));   // src/ram.vhd(56[12:17])
    SB_DFF i6017_6018 (.Q(ram_s_250_1), .C(CLK_3P3_MHZ_c), .D(n2889));   // src/ram.vhd(56[12:17])
    SB_DFF i6014_6015 (.Q(ram_s_250_0), .C(CLK_3P3_MHZ_c), .D(n2888));   // src/ram.vhd(56[12:17])
    SB_DFF i6011_6012 (.Q(ram_s_249_7), .C(CLK_3P3_MHZ_c), .D(n2887));   // src/ram.vhd(56[12:17])
    SB_DFF i6008_6009 (.Q(ram_s_249_6), .C(CLK_3P3_MHZ_c), .D(n2886));   // src/ram.vhd(56[12:17])
    SB_DFF i6005_6006 (.Q(ram_s_249_5), .C(CLK_3P3_MHZ_c), .D(n2885));   // src/ram.vhd(56[12:17])
    SB_DFF i6002_6003 (.Q(ram_s_249_4), .C(CLK_3P3_MHZ_c), .D(n2884));   // src/ram.vhd(56[12:17])
    SB_DFF i5999_6000 (.Q(ram_s_249_3), .C(CLK_3P3_MHZ_c), .D(n2883));   // src/ram.vhd(56[12:17])
    SB_DFF i5996_5997 (.Q(ram_s_249_2), .C(CLK_3P3_MHZ_c), .D(n2882));   // src/ram.vhd(56[12:17])
    SB_DFF i5993_5994 (.Q(ram_s_249_1), .C(CLK_3P3_MHZ_c), .D(n2881));   // src/ram.vhd(56[12:17])
    SB_DFF i5990_5991 (.Q(ram_s_249_0), .C(CLK_3P3_MHZ_c), .D(n2880));   // src/ram.vhd(56[12:17])
    SB_DFF i5987_5988 (.Q(ram_s_248_7), .C(CLK_3P3_MHZ_c), .D(n2879));   // src/ram.vhd(56[12:17])
    SB_DFF i5984_5985 (.Q(ram_s_248_6), .C(CLK_3P3_MHZ_c), .D(n2878));   // src/ram.vhd(56[12:17])
    SB_DFF i5981_5982 (.Q(ram_s_248_5), .C(CLK_3P3_MHZ_c), .D(n2877));   // src/ram.vhd(56[12:17])
    SB_DFF i5978_5979 (.Q(ram_s_248_4), .C(CLK_3P3_MHZ_c), .D(n2876));   // src/ram.vhd(56[12:17])
    SB_DFF i5975_5976 (.Q(ram_s_248_3), .C(CLK_3P3_MHZ_c), .D(n2875));   // src/ram.vhd(56[12:17])
    SB_DFF i5972_5973 (.Q(ram_s_248_2), .C(CLK_3P3_MHZ_c), .D(n2874));   // src/ram.vhd(56[12:17])
    SB_DFF i5969_5970 (.Q(ram_s_248_1), .C(CLK_3P3_MHZ_c), .D(n2873));   // src/ram.vhd(56[12:17])
    SB_DFF i5966_5967 (.Q(ram_s_248_0), .C(CLK_3P3_MHZ_c), .D(n2872));   // src/ram.vhd(56[12:17])
    SB_DFF i5963_5964 (.Q(ram_s_247_7), .C(CLK_3P3_MHZ_c), .D(n2871));   // src/ram.vhd(56[12:17])
    SB_DFF i5960_5961 (.Q(ram_s_247_6), .C(CLK_3P3_MHZ_c), .D(n2870));   // src/ram.vhd(56[12:17])
    SB_DFF i5957_5958 (.Q(ram_s_247_5), .C(CLK_3P3_MHZ_c), .D(n2869));   // src/ram.vhd(56[12:17])
    SB_DFF i5954_5955 (.Q(ram_s_247_4), .C(CLK_3P3_MHZ_c), .D(n2868));   // src/ram.vhd(56[12:17])
    SB_DFF i5951_5952 (.Q(ram_s_247_3), .C(CLK_3P3_MHZ_c), .D(n2867));   // src/ram.vhd(56[12:17])
    SB_DFF i5948_5949 (.Q(ram_s_247_2), .C(CLK_3P3_MHZ_c), .D(n2866));   // src/ram.vhd(56[12:17])
    SB_DFF i5945_5946 (.Q(ram_s_247_1), .C(CLK_3P3_MHZ_c), .D(n2865));   // src/ram.vhd(56[12:17])
    SB_DFF i5942_5943 (.Q(ram_s_247_0), .C(CLK_3P3_MHZ_c), .D(n2864));   // src/ram.vhd(56[12:17])
    SB_DFF i5939_5940 (.Q(ram_s_246_7), .C(CLK_3P3_MHZ_c), .D(n2863));   // src/ram.vhd(56[12:17])
    SB_DFF i5936_5937 (.Q(ram_s_246_6), .C(CLK_3P3_MHZ_c), .D(n2862));   // src/ram.vhd(56[12:17])
    SB_DFF i5933_5934 (.Q(ram_s_246_5), .C(CLK_3P3_MHZ_c), .D(n2861));   // src/ram.vhd(56[12:17])
    SB_DFF i5930_5931 (.Q(ram_s_246_4), .C(CLK_3P3_MHZ_c), .D(n2860));   // src/ram.vhd(56[12:17])
    SB_DFF i5927_5928 (.Q(ram_s_246_3), .C(CLK_3P3_MHZ_c), .D(n2859));   // src/ram.vhd(56[12:17])
    SB_DFF i5924_5925 (.Q(ram_s_246_2), .C(CLK_3P3_MHZ_c), .D(n2858));   // src/ram.vhd(56[12:17])
    SB_DFF i5921_5922 (.Q(ram_s_246_1), .C(CLK_3P3_MHZ_c), .D(n2857));   // src/ram.vhd(56[12:17])
    SB_DFF i5918_5919 (.Q(ram_s_246_0), .C(CLK_3P3_MHZ_c), .D(n2856));   // src/ram.vhd(56[12:17])
    SB_DFF i5915_5916 (.Q(ram_s_245_7), .C(CLK_3P3_MHZ_c), .D(n2855));   // src/ram.vhd(56[12:17])
    SB_DFF i5912_5913 (.Q(ram_s_245_6), .C(CLK_3P3_MHZ_c), .D(n2854));   // src/ram.vhd(56[12:17])
    SB_DFF i5909_5910 (.Q(ram_s_245_5), .C(CLK_3P3_MHZ_c), .D(n2853));   // src/ram.vhd(56[12:17])
    SB_DFF i5906_5907 (.Q(ram_s_245_4), .C(CLK_3P3_MHZ_c), .D(n2852));   // src/ram.vhd(56[12:17])
    SB_DFF i5903_5904 (.Q(ram_s_245_3), .C(CLK_3P3_MHZ_c), .D(n2851));   // src/ram.vhd(56[12:17])
    SB_DFF i5900_5901 (.Q(ram_s_245_2), .C(CLK_3P3_MHZ_c), .D(n2850));   // src/ram.vhd(56[12:17])
    SB_DFF i5897_5898 (.Q(ram_s_245_1), .C(CLK_3P3_MHZ_c), .D(n2849));   // src/ram.vhd(56[12:17])
    SB_DFF i5894_5895 (.Q(ram_s_245_0), .C(CLK_3P3_MHZ_c), .D(n2848));   // src/ram.vhd(56[12:17])
    SB_DFF i5891_5892 (.Q(ram_s_244_7), .C(CLK_3P3_MHZ_c), .D(n2847));   // src/ram.vhd(56[12:17])
    SB_DFF i5888_5889 (.Q(ram_s_244_6), .C(CLK_3P3_MHZ_c), .D(n2846));   // src/ram.vhd(56[12:17])
    SB_DFF i5885_5886 (.Q(ram_s_244_5), .C(CLK_3P3_MHZ_c), .D(n2845));   // src/ram.vhd(56[12:17])
    SB_DFF i5882_5883 (.Q(ram_s_244_4), .C(CLK_3P3_MHZ_c), .D(n2844));   // src/ram.vhd(56[12:17])
    SB_DFF i5879_5880 (.Q(ram_s_244_3), .C(CLK_3P3_MHZ_c), .D(n2843));   // src/ram.vhd(56[12:17])
    SB_DFF i5876_5877 (.Q(ram_s_244_2), .C(CLK_3P3_MHZ_c), .D(n2842));   // src/ram.vhd(56[12:17])
    SB_DFF i5873_5874 (.Q(ram_s_244_1), .C(CLK_3P3_MHZ_c), .D(n2841));   // src/ram.vhd(56[12:17])
    SB_DFF i5870_5871 (.Q(ram_s_244_0), .C(CLK_3P3_MHZ_c), .D(n2840));   // src/ram.vhd(56[12:17])
    SB_DFF i5867_5868 (.Q(ram_s_243_7), .C(CLK_3P3_MHZ_c), .D(n2839));   // src/ram.vhd(56[12:17])
    SB_DFF i5864_5865 (.Q(ram_s_243_6), .C(CLK_3P3_MHZ_c), .D(n2838));   // src/ram.vhd(56[12:17])
    SB_DFF i5861_5862 (.Q(ram_s_243_5), .C(CLK_3P3_MHZ_c), .D(n2837));   // src/ram.vhd(56[12:17])
    SB_DFF i5858_5859 (.Q(ram_s_243_4), .C(CLK_3P3_MHZ_c), .D(n2836));   // src/ram.vhd(56[12:17])
    SB_DFF i5855_5856 (.Q(ram_s_243_3), .C(CLK_3P3_MHZ_c), .D(n2835));   // src/ram.vhd(56[12:17])
    SB_DFF i5852_5853 (.Q(ram_s_243_2), .C(CLK_3P3_MHZ_c), .D(n2834));   // src/ram.vhd(56[12:17])
    SB_DFF i5849_5850 (.Q(ram_s_243_1), .C(CLK_3P3_MHZ_c), .D(n2833));   // src/ram.vhd(56[12:17])
    SB_DFF i5846_5847 (.Q(ram_s_243_0), .C(CLK_3P3_MHZ_c), .D(n2832));   // src/ram.vhd(56[12:17])
    SB_DFF i5843_5844 (.Q(ram_s_242_7), .C(CLK_3P3_MHZ_c), .D(n2831));   // src/ram.vhd(56[12:17])
    SB_DFF i5840_5841 (.Q(ram_s_242_6), .C(CLK_3P3_MHZ_c), .D(n2830));   // src/ram.vhd(56[12:17])
    SB_DFF i5837_5838 (.Q(ram_s_242_5), .C(CLK_3P3_MHZ_c), .D(n2829));   // src/ram.vhd(56[12:17])
    SB_DFF i5834_5835 (.Q(ram_s_242_4), .C(CLK_3P3_MHZ_c), .D(n2828));   // src/ram.vhd(56[12:17])
    SB_DFF i5831_5832 (.Q(ram_s_242_3), .C(CLK_3P3_MHZ_c), .D(n2827));   // src/ram.vhd(56[12:17])
    SB_DFF i5828_5829 (.Q(ram_s_242_2), .C(CLK_3P3_MHZ_c), .D(n2826));   // src/ram.vhd(56[12:17])
    SB_DFF i5825_5826 (.Q(ram_s_242_1), .C(CLK_3P3_MHZ_c), .D(n2825));   // src/ram.vhd(56[12:17])
    SB_DFF i5822_5823 (.Q(ram_s_242_0), .C(CLK_3P3_MHZ_c), .D(n2824));   // src/ram.vhd(56[12:17])
    SB_DFF i5819_5820 (.Q(ram_s_241_7), .C(CLK_3P3_MHZ_c), .D(n2823));   // src/ram.vhd(56[12:17])
    SB_DFF i5816_5817 (.Q(ram_s_241_6), .C(CLK_3P3_MHZ_c), .D(n2822));   // src/ram.vhd(56[12:17])
    SB_DFF i5813_5814 (.Q(ram_s_241_5), .C(CLK_3P3_MHZ_c), .D(n2821));   // src/ram.vhd(56[12:17])
    SB_DFF i5810_5811 (.Q(ram_s_241_4), .C(CLK_3P3_MHZ_c), .D(n2820));   // src/ram.vhd(56[12:17])
    SB_DFF i5807_5808 (.Q(ram_s_241_3), .C(CLK_3P3_MHZ_c), .D(n2819));   // src/ram.vhd(56[12:17])
    SB_DFF i5804_5805 (.Q(ram_s_241_2), .C(CLK_3P3_MHZ_c), .D(n2818));   // src/ram.vhd(56[12:17])
    SB_DFF i5801_5802 (.Q(ram_s_241_1), .C(CLK_3P3_MHZ_c), .D(n2817));   // src/ram.vhd(56[12:17])
    SB_DFF i5798_5799 (.Q(ram_s_241_0), .C(CLK_3P3_MHZ_c), .D(n2816));   // src/ram.vhd(56[12:17])
    SB_DFF i5795_5796 (.Q(ram_s_240_7), .C(CLK_3P3_MHZ_c), .D(n2815));   // src/ram.vhd(56[12:17])
    SB_DFF i5792_5793 (.Q(ram_s_240_6), .C(CLK_3P3_MHZ_c), .D(n2814));   // src/ram.vhd(56[12:17])
    SB_DFF i5789_5790 (.Q(ram_s_240_5), .C(CLK_3P3_MHZ_c), .D(n2813));   // src/ram.vhd(56[12:17])
    SB_DFF i5786_5787 (.Q(ram_s_240_4), .C(CLK_3P3_MHZ_c), .D(n2812));   // src/ram.vhd(56[12:17])
    SB_DFF i5783_5784 (.Q(ram_s_240_3), .C(CLK_3P3_MHZ_c), .D(n2811));   // src/ram.vhd(56[12:17])
    SB_DFF i5780_5781 (.Q(ram_s_240_2), .C(CLK_3P3_MHZ_c), .D(n2810));   // src/ram.vhd(56[12:17])
    SB_DFF i5777_5778 (.Q(ram_s_240_1), .C(CLK_3P3_MHZ_c), .D(n2809));   // src/ram.vhd(56[12:17])
    SB_DFF i5774_5775 (.Q(ram_s_240_0), .C(CLK_3P3_MHZ_c), .D(n2808));   // src/ram.vhd(56[12:17])
    SB_DFF i5771_5772 (.Q(ram_s_239_7), .C(CLK_3P3_MHZ_c), .D(n2807));   // src/ram.vhd(56[12:17])
    SB_DFF i5768_5769 (.Q(ram_s_239_6), .C(CLK_3P3_MHZ_c), .D(n2806));   // src/ram.vhd(56[12:17])
    SB_DFF i5765_5766 (.Q(ram_s_239_5), .C(CLK_3P3_MHZ_c), .D(n2805));   // src/ram.vhd(56[12:17])
    SB_DFF i5762_5763 (.Q(ram_s_239_4), .C(CLK_3P3_MHZ_c), .D(n2804));   // src/ram.vhd(56[12:17])
    SB_DFF i5759_5760 (.Q(ram_s_239_3), .C(CLK_3P3_MHZ_c), .D(n2803));   // src/ram.vhd(56[12:17])
    SB_DFF i5756_5757 (.Q(ram_s_239_2), .C(CLK_3P3_MHZ_c), .D(n2802));   // src/ram.vhd(56[12:17])
    SB_DFF i5753_5754 (.Q(ram_s_239_1), .C(CLK_3P3_MHZ_c), .D(n2801));   // src/ram.vhd(56[12:17])
    SB_DFF i5750_5751 (.Q(ram_s_239_0), .C(CLK_3P3_MHZ_c), .D(n2800));   // src/ram.vhd(56[12:17])
    SB_DFF i5747_5748 (.Q(ram_s_238_7), .C(CLK_3P3_MHZ_c), .D(n2799));   // src/ram.vhd(56[12:17])
    SB_DFF i5744_5745 (.Q(ram_s_238_6), .C(CLK_3P3_MHZ_c), .D(n2798));   // src/ram.vhd(56[12:17])
    SB_DFF i5741_5742 (.Q(ram_s_238_5), .C(CLK_3P3_MHZ_c), .D(n2797));   // src/ram.vhd(56[12:17])
    SB_DFF i5738_5739 (.Q(ram_s_238_4), .C(CLK_3P3_MHZ_c), .D(n2796));   // src/ram.vhd(56[12:17])
    SB_DFF i5735_5736 (.Q(ram_s_238_3), .C(CLK_3P3_MHZ_c), .D(n2795));   // src/ram.vhd(56[12:17])
    SB_DFF i5732_5733 (.Q(ram_s_238_2), .C(CLK_3P3_MHZ_c), .D(n2794));   // src/ram.vhd(56[12:17])
    SB_DFF i5729_5730 (.Q(ram_s_238_1), .C(CLK_3P3_MHZ_c), .D(n2793));   // src/ram.vhd(56[12:17])
    SB_DFF i5726_5727 (.Q(ram_s_238_0), .C(CLK_3P3_MHZ_c), .D(n2792));   // src/ram.vhd(56[12:17])
    SB_DFF i5723_5724 (.Q(ram_s_237_7), .C(CLK_3P3_MHZ_c), .D(n2791));   // src/ram.vhd(56[12:17])
    SB_DFF i5720_5721 (.Q(ram_s_237_6), .C(CLK_3P3_MHZ_c), .D(n2790));   // src/ram.vhd(56[12:17])
    SB_DFF i5717_5718 (.Q(ram_s_237_5), .C(CLK_3P3_MHZ_c), .D(n2789));   // src/ram.vhd(56[12:17])
    SB_DFF i5714_5715 (.Q(ram_s_237_4), .C(CLK_3P3_MHZ_c), .D(n2788));   // src/ram.vhd(56[12:17])
    SB_DFF i5711_5712 (.Q(ram_s_237_3), .C(CLK_3P3_MHZ_c), .D(n2787));   // src/ram.vhd(56[12:17])
    SB_DFF i5708_5709 (.Q(ram_s_237_2), .C(CLK_3P3_MHZ_c), .D(n2786));   // src/ram.vhd(56[12:17])
    SB_DFF i5705_5706 (.Q(ram_s_237_1), .C(CLK_3P3_MHZ_c), .D(n2785));   // src/ram.vhd(56[12:17])
    SB_DFF i5702_5703 (.Q(ram_s_237_0), .C(CLK_3P3_MHZ_c), .D(n2784));   // src/ram.vhd(56[12:17])
    SB_DFF i5699_5700 (.Q(ram_s_236_7), .C(CLK_3P3_MHZ_c), .D(n2783));   // src/ram.vhd(56[12:17])
    SB_DFF i5696_5697 (.Q(ram_s_236_6), .C(CLK_3P3_MHZ_c), .D(n2782));   // src/ram.vhd(56[12:17])
    SB_DFF i5693_5694 (.Q(ram_s_236_5), .C(CLK_3P3_MHZ_c), .D(n2781));   // src/ram.vhd(56[12:17])
    SB_DFF i5690_5691 (.Q(ram_s_236_4), .C(CLK_3P3_MHZ_c), .D(n2780));   // src/ram.vhd(56[12:17])
    SB_DFF i5687_5688 (.Q(ram_s_236_3), .C(CLK_3P3_MHZ_c), .D(n2779));   // src/ram.vhd(56[12:17])
    SB_DFF i5684_5685 (.Q(ram_s_236_2), .C(CLK_3P3_MHZ_c), .D(n2778));   // src/ram.vhd(56[12:17])
    SB_DFF i5681_5682 (.Q(ram_s_236_1), .C(CLK_3P3_MHZ_c), .D(n2777));   // src/ram.vhd(56[12:17])
    SB_DFF i5678_5679 (.Q(ram_s_236_0), .C(CLK_3P3_MHZ_c), .D(n2776));   // src/ram.vhd(56[12:17])
    SB_DFF i5675_5676 (.Q(ram_s_235_7), .C(CLK_3P3_MHZ_c), .D(n2775));   // src/ram.vhd(56[12:17])
    SB_DFF i5672_5673 (.Q(ram_s_235_6), .C(CLK_3P3_MHZ_c), .D(n2774));   // src/ram.vhd(56[12:17])
    SB_DFF i5669_5670 (.Q(ram_s_235_5), .C(CLK_3P3_MHZ_c), .D(n2773));   // src/ram.vhd(56[12:17])
    SB_DFF i5666_5667 (.Q(ram_s_235_4), .C(CLK_3P3_MHZ_c), .D(n2772));   // src/ram.vhd(56[12:17])
    SB_DFF i5663_5664 (.Q(ram_s_235_3), .C(CLK_3P3_MHZ_c), .D(n2771));   // src/ram.vhd(56[12:17])
    SB_DFF i5660_5661 (.Q(ram_s_235_2), .C(CLK_3P3_MHZ_c), .D(n2770));   // src/ram.vhd(56[12:17])
    SB_DFF i5657_5658 (.Q(ram_s_235_1), .C(CLK_3P3_MHZ_c), .D(n2769));   // src/ram.vhd(56[12:17])
    SB_DFF i5654_5655 (.Q(ram_s_235_0), .C(CLK_3P3_MHZ_c), .D(n2768));   // src/ram.vhd(56[12:17])
    SB_DFF i5651_5652 (.Q(ram_s_234_7), .C(CLK_3P3_MHZ_c), .D(n2767));   // src/ram.vhd(56[12:17])
    SB_DFF i5648_5649 (.Q(ram_s_234_6), .C(CLK_3P3_MHZ_c), .D(n2766));   // src/ram.vhd(56[12:17])
    SB_DFF i5645_5646 (.Q(ram_s_234_5), .C(CLK_3P3_MHZ_c), .D(n2765));   // src/ram.vhd(56[12:17])
    SB_DFF i5642_5643 (.Q(ram_s_234_4), .C(CLK_3P3_MHZ_c), .D(n2764));   // src/ram.vhd(56[12:17])
    SB_DFF i5639_5640 (.Q(ram_s_234_3), .C(CLK_3P3_MHZ_c), .D(n2763));   // src/ram.vhd(56[12:17])
    SB_DFF i5636_5637 (.Q(ram_s_234_2), .C(CLK_3P3_MHZ_c), .D(n2762));   // src/ram.vhd(56[12:17])
    SB_DFF i5633_5634 (.Q(ram_s_234_1), .C(CLK_3P3_MHZ_c), .D(n2761));   // src/ram.vhd(56[12:17])
    SB_DFF i5630_5631 (.Q(ram_s_234_0), .C(CLK_3P3_MHZ_c), .D(n2760));   // src/ram.vhd(56[12:17])
    SB_DFF i5627_5628 (.Q(ram_s_233_7), .C(CLK_3P3_MHZ_c), .D(n2759));   // src/ram.vhd(56[12:17])
    SB_DFF i5624_5625 (.Q(ram_s_233_6), .C(CLK_3P3_MHZ_c), .D(n2758));   // src/ram.vhd(56[12:17])
    SB_DFF i5621_5622 (.Q(ram_s_233_5), .C(CLK_3P3_MHZ_c), .D(n2757));   // src/ram.vhd(56[12:17])
    SB_DFF i5618_5619 (.Q(ram_s_233_4), .C(CLK_3P3_MHZ_c), .D(n2756));   // src/ram.vhd(56[12:17])
    SB_DFF i5615_5616 (.Q(ram_s_233_3), .C(CLK_3P3_MHZ_c), .D(n2755));   // src/ram.vhd(56[12:17])
    SB_DFF i5612_5613 (.Q(ram_s_233_2), .C(CLK_3P3_MHZ_c), .D(n2754));   // src/ram.vhd(56[12:17])
    SB_DFF i5609_5610 (.Q(ram_s_233_1), .C(CLK_3P3_MHZ_c), .D(n2753));   // src/ram.vhd(56[12:17])
    SB_DFF i5606_5607 (.Q(ram_s_233_0), .C(CLK_3P3_MHZ_c), .D(n2752));   // src/ram.vhd(56[12:17])
    SB_DFF i5603_5604 (.Q(ram_s_232_7), .C(CLK_3P3_MHZ_c), .D(n2751));   // src/ram.vhd(56[12:17])
    SB_DFF i5600_5601 (.Q(ram_s_232_6), .C(CLK_3P3_MHZ_c), .D(n2750));   // src/ram.vhd(56[12:17])
    SB_DFF i5597_5598 (.Q(ram_s_232_5), .C(CLK_3P3_MHZ_c), .D(n2749));   // src/ram.vhd(56[12:17])
    SB_DFF i5594_5595 (.Q(ram_s_232_4), .C(CLK_3P3_MHZ_c), .D(n2748));   // src/ram.vhd(56[12:17])
    SB_DFF i5591_5592 (.Q(ram_s_232_3), .C(CLK_3P3_MHZ_c), .D(n2747));   // src/ram.vhd(56[12:17])
    SB_DFF i5588_5589 (.Q(ram_s_232_2), .C(CLK_3P3_MHZ_c), .D(n2746));   // src/ram.vhd(56[12:17])
    SB_DFF i5585_5586 (.Q(ram_s_232_1), .C(CLK_3P3_MHZ_c), .D(n2745));   // src/ram.vhd(56[12:17])
    SB_DFF i5582_5583 (.Q(ram_s_232_0), .C(CLK_3P3_MHZ_c), .D(n2744));   // src/ram.vhd(56[12:17])
    SB_DFF i5579_5580 (.Q(ram_s_231_7), .C(CLK_3P3_MHZ_c), .D(n2743));   // src/ram.vhd(56[12:17])
    SB_DFF i5576_5577 (.Q(ram_s_231_6), .C(CLK_3P3_MHZ_c), .D(n2742));   // src/ram.vhd(56[12:17])
    SB_DFF i5573_5574 (.Q(ram_s_231_5), .C(CLK_3P3_MHZ_c), .D(n2741));   // src/ram.vhd(56[12:17])
    SB_DFF i5570_5571 (.Q(ram_s_231_4), .C(CLK_3P3_MHZ_c), .D(n2740));   // src/ram.vhd(56[12:17])
    SB_DFF i5567_5568 (.Q(ram_s_231_3), .C(CLK_3P3_MHZ_c), .D(n2739));   // src/ram.vhd(56[12:17])
    SB_DFF i5564_5565 (.Q(ram_s_231_2), .C(CLK_3P3_MHZ_c), .D(n2738));   // src/ram.vhd(56[12:17])
    SB_DFF i5561_5562 (.Q(ram_s_231_1), .C(CLK_3P3_MHZ_c), .D(n2737));   // src/ram.vhd(56[12:17])
    SB_DFF i5558_5559 (.Q(ram_s_231_0), .C(CLK_3P3_MHZ_c), .D(n2736));   // src/ram.vhd(56[12:17])
    SB_DFF i5555_5556 (.Q(ram_s_230_7), .C(CLK_3P3_MHZ_c), .D(n2735));   // src/ram.vhd(56[12:17])
    SB_DFF i5552_5553 (.Q(ram_s_230_6), .C(CLK_3P3_MHZ_c), .D(n2734));   // src/ram.vhd(56[12:17])
    SB_DFF i5549_5550 (.Q(ram_s_230_5), .C(CLK_3P3_MHZ_c), .D(n2733));   // src/ram.vhd(56[12:17])
    SB_DFF i5546_5547 (.Q(ram_s_230_4), .C(CLK_3P3_MHZ_c), .D(n2732));   // src/ram.vhd(56[12:17])
    SB_DFF i5543_5544 (.Q(ram_s_230_3), .C(CLK_3P3_MHZ_c), .D(n2731));   // src/ram.vhd(56[12:17])
    SB_DFF i5540_5541 (.Q(ram_s_230_2), .C(CLK_3P3_MHZ_c), .D(n2730));   // src/ram.vhd(56[12:17])
    SB_DFF i5537_5538 (.Q(ram_s_230_1), .C(CLK_3P3_MHZ_c), .D(n2729));   // src/ram.vhd(56[12:17])
    SB_DFF i5534_5535 (.Q(ram_s_230_0), .C(CLK_3P3_MHZ_c), .D(n2728));   // src/ram.vhd(56[12:17])
    SB_DFF i5531_5532 (.Q(ram_s_229_7), .C(CLK_3P3_MHZ_c), .D(n2727));   // src/ram.vhd(56[12:17])
    SB_DFF i5528_5529 (.Q(ram_s_229_6), .C(CLK_3P3_MHZ_c), .D(n2726));   // src/ram.vhd(56[12:17])
    SB_DFF i5525_5526 (.Q(ram_s_229_5), .C(CLK_3P3_MHZ_c), .D(n2725));   // src/ram.vhd(56[12:17])
    SB_DFF i5522_5523 (.Q(ram_s_229_4), .C(CLK_3P3_MHZ_c), .D(n2724));   // src/ram.vhd(56[12:17])
    SB_DFF i5519_5520 (.Q(ram_s_229_3), .C(CLK_3P3_MHZ_c), .D(n2723));   // src/ram.vhd(56[12:17])
    SB_DFF i5516_5517 (.Q(ram_s_229_2), .C(CLK_3P3_MHZ_c), .D(n2722));   // src/ram.vhd(56[12:17])
    SB_DFF i5513_5514 (.Q(ram_s_229_1), .C(CLK_3P3_MHZ_c), .D(n2721));   // src/ram.vhd(56[12:17])
    SB_DFF i5510_5511 (.Q(ram_s_229_0), .C(CLK_3P3_MHZ_c), .D(n2720));   // src/ram.vhd(56[12:17])
    SB_DFF i5507_5508 (.Q(ram_s_228_7), .C(CLK_3P3_MHZ_c), .D(n2719));   // src/ram.vhd(56[12:17])
    SB_DFF i5504_5505 (.Q(ram_s_228_6), .C(CLK_3P3_MHZ_c), .D(n2718));   // src/ram.vhd(56[12:17])
    SB_DFF i5501_5502 (.Q(ram_s_228_5), .C(CLK_3P3_MHZ_c), .D(n2717));   // src/ram.vhd(56[12:17])
    SB_DFF i5498_5499 (.Q(ram_s_228_4), .C(CLK_3P3_MHZ_c), .D(n2716));   // src/ram.vhd(56[12:17])
    SB_DFF i5495_5496 (.Q(ram_s_228_3), .C(CLK_3P3_MHZ_c), .D(n2715));   // src/ram.vhd(56[12:17])
    SB_DFF i5492_5493 (.Q(ram_s_228_2), .C(CLK_3P3_MHZ_c), .D(n2714));   // src/ram.vhd(56[12:17])
    SB_DFF i5489_5490 (.Q(ram_s_228_1), .C(CLK_3P3_MHZ_c), .D(n2713));   // src/ram.vhd(56[12:17])
    SB_DFF i5486_5487 (.Q(ram_s_228_0), .C(CLK_3P3_MHZ_c), .D(n2712));   // src/ram.vhd(56[12:17])
    SB_DFF i5483_5484 (.Q(ram_s_227_7), .C(CLK_3P3_MHZ_c), .D(n2711));   // src/ram.vhd(56[12:17])
    SB_DFF i5480_5481 (.Q(ram_s_227_6), .C(CLK_3P3_MHZ_c), .D(n2710));   // src/ram.vhd(56[12:17])
    SB_DFF i5477_5478 (.Q(ram_s_227_5), .C(CLK_3P3_MHZ_c), .D(n2709));   // src/ram.vhd(56[12:17])
    SB_DFF i5474_5475 (.Q(ram_s_227_4), .C(CLK_3P3_MHZ_c), .D(n2708));   // src/ram.vhd(56[12:17])
    SB_DFF i5471_5472 (.Q(ram_s_227_3), .C(CLK_3P3_MHZ_c), .D(n2707));   // src/ram.vhd(56[12:17])
    SB_DFF i5468_5469 (.Q(ram_s_227_2), .C(CLK_3P3_MHZ_c), .D(n2706));   // src/ram.vhd(56[12:17])
    SB_DFF i5465_5466 (.Q(ram_s_227_1), .C(CLK_3P3_MHZ_c), .D(n2705));   // src/ram.vhd(56[12:17])
    SB_DFF i5462_5463 (.Q(ram_s_227_0), .C(CLK_3P3_MHZ_c), .D(n2704));   // src/ram.vhd(56[12:17])
    SB_DFF i5459_5460 (.Q(ram_s_226_7), .C(CLK_3P3_MHZ_c), .D(n2703));   // src/ram.vhd(56[12:17])
    SB_DFF i5456_5457 (.Q(ram_s_226_6), .C(CLK_3P3_MHZ_c), .D(n2702));   // src/ram.vhd(56[12:17])
    SB_DFF i5453_5454 (.Q(ram_s_226_5), .C(CLK_3P3_MHZ_c), .D(n2701));   // src/ram.vhd(56[12:17])
    SB_DFF i5450_5451 (.Q(ram_s_226_4), .C(CLK_3P3_MHZ_c), .D(n2700));   // src/ram.vhd(56[12:17])
    SB_DFF i5447_5448 (.Q(ram_s_226_3), .C(CLK_3P3_MHZ_c), .D(n2699));   // src/ram.vhd(56[12:17])
    SB_DFF i5444_5445 (.Q(ram_s_226_2), .C(CLK_3P3_MHZ_c), .D(n2698));   // src/ram.vhd(56[12:17])
    SB_DFF i5441_5442 (.Q(ram_s_226_1), .C(CLK_3P3_MHZ_c), .D(n2697));   // src/ram.vhd(56[12:17])
    SB_DFF i5438_5439 (.Q(ram_s_226_0), .C(CLK_3P3_MHZ_c), .D(n2696));   // src/ram.vhd(56[12:17])
    SB_DFF i5435_5436 (.Q(ram_s_225_7), .C(CLK_3P3_MHZ_c), .D(n2695));   // src/ram.vhd(56[12:17])
    SB_DFF i5432_5433 (.Q(ram_s_225_6), .C(CLK_3P3_MHZ_c), .D(n2694));   // src/ram.vhd(56[12:17])
    SB_DFF i5429_5430 (.Q(ram_s_225_5), .C(CLK_3P3_MHZ_c), .D(n2693));   // src/ram.vhd(56[12:17])
    SB_DFF i5426_5427 (.Q(ram_s_225_4), .C(CLK_3P3_MHZ_c), .D(n2692));   // src/ram.vhd(56[12:17])
    SB_DFF i5423_5424 (.Q(ram_s_225_3), .C(CLK_3P3_MHZ_c), .D(n2691));   // src/ram.vhd(56[12:17])
    SB_DFF i5420_5421 (.Q(ram_s_225_2), .C(CLK_3P3_MHZ_c), .D(n2690));   // src/ram.vhd(56[12:17])
    SB_DFF i5417_5418 (.Q(ram_s_225_1), .C(CLK_3P3_MHZ_c), .D(n2689));   // src/ram.vhd(56[12:17])
    SB_DFF i5414_5415 (.Q(ram_s_225_0), .C(CLK_3P3_MHZ_c), .D(n2688));   // src/ram.vhd(56[12:17])
    SB_DFF i5411_5412 (.Q(ram_s_224_7), .C(CLK_3P3_MHZ_c), .D(n2687));   // src/ram.vhd(56[12:17])
    SB_DFF i5408_5409 (.Q(ram_s_224_6), .C(CLK_3P3_MHZ_c), .D(n2686));   // src/ram.vhd(56[12:17])
    SB_DFF i5405_5406 (.Q(ram_s_224_5), .C(CLK_3P3_MHZ_c), .D(n2685));   // src/ram.vhd(56[12:17])
    SB_DFF i5402_5403 (.Q(ram_s_224_4), .C(CLK_3P3_MHZ_c), .D(n2684));   // src/ram.vhd(56[12:17])
    SB_DFF i5399_5400 (.Q(ram_s_224_3), .C(CLK_3P3_MHZ_c), .D(n2683));   // src/ram.vhd(56[12:17])
    SB_DFF i5396_5397 (.Q(ram_s_224_2), .C(CLK_3P3_MHZ_c), .D(n2682));   // src/ram.vhd(56[12:17])
    SB_DFF i5393_5394 (.Q(ram_s_224_1), .C(CLK_3P3_MHZ_c), .D(n2681));   // src/ram.vhd(56[12:17])
    SB_DFF i5390_5391 (.Q(ram_s_224_0), .C(CLK_3P3_MHZ_c), .D(n2680));   // src/ram.vhd(56[12:17])
    SB_DFF i5387_5388 (.Q(ram_s_223_7), .C(CLK_3P3_MHZ_c), .D(n2679));   // src/ram.vhd(56[12:17])
    SB_DFF i5384_5385 (.Q(ram_s_223_6), .C(CLK_3P3_MHZ_c), .D(n2678));   // src/ram.vhd(56[12:17])
    SB_DFF i5381_5382 (.Q(ram_s_223_5), .C(CLK_3P3_MHZ_c), .D(n2677));   // src/ram.vhd(56[12:17])
    SB_DFF i5378_5379 (.Q(ram_s_223_4), .C(CLK_3P3_MHZ_c), .D(n2676));   // src/ram.vhd(56[12:17])
    SB_DFF i5375_5376 (.Q(ram_s_223_3), .C(CLK_3P3_MHZ_c), .D(n2675));   // src/ram.vhd(56[12:17])
    SB_DFF i5372_5373 (.Q(ram_s_223_2), .C(CLK_3P3_MHZ_c), .D(n2674));   // src/ram.vhd(56[12:17])
    SB_DFF i5369_5370 (.Q(ram_s_223_1), .C(CLK_3P3_MHZ_c), .D(n2673));   // src/ram.vhd(56[12:17])
    SB_DFF i5366_5367 (.Q(ram_s_223_0), .C(CLK_3P3_MHZ_c), .D(n2672));   // src/ram.vhd(56[12:17])
    SB_DFF i5363_5364 (.Q(ram_s_222_7), .C(CLK_3P3_MHZ_c), .D(n2671));   // src/ram.vhd(56[12:17])
    SB_DFF i5360_5361 (.Q(ram_s_222_6), .C(CLK_3P3_MHZ_c), .D(n2670));   // src/ram.vhd(56[12:17])
    SB_DFF i5357_5358 (.Q(ram_s_222_5), .C(CLK_3P3_MHZ_c), .D(n2669));   // src/ram.vhd(56[12:17])
    SB_DFF i5354_5355 (.Q(ram_s_222_4), .C(CLK_3P3_MHZ_c), .D(n2668));   // src/ram.vhd(56[12:17])
    SB_DFF i5351_5352 (.Q(ram_s_222_3), .C(CLK_3P3_MHZ_c), .D(n2667));   // src/ram.vhd(56[12:17])
    SB_DFF i5348_5349 (.Q(ram_s_222_2), .C(CLK_3P3_MHZ_c), .D(n2666));   // src/ram.vhd(56[12:17])
    SB_DFF i5345_5346 (.Q(ram_s_222_1), .C(CLK_3P3_MHZ_c), .D(n2665));   // src/ram.vhd(56[12:17])
    SB_DFF i5342_5343 (.Q(ram_s_222_0), .C(CLK_3P3_MHZ_c), .D(n2664));   // src/ram.vhd(56[12:17])
    SB_DFF i5339_5340 (.Q(ram_s_221_7), .C(CLK_3P3_MHZ_c), .D(n2663));   // src/ram.vhd(56[12:17])
    SB_DFF i5336_5337 (.Q(ram_s_221_6), .C(CLK_3P3_MHZ_c), .D(n2662));   // src/ram.vhd(56[12:17])
    SB_DFF i5333_5334 (.Q(ram_s_221_5), .C(CLK_3P3_MHZ_c), .D(n2661));   // src/ram.vhd(56[12:17])
    SB_DFF i5330_5331 (.Q(ram_s_221_4), .C(CLK_3P3_MHZ_c), .D(n2660));   // src/ram.vhd(56[12:17])
    SB_DFF i5327_5328 (.Q(ram_s_221_3), .C(CLK_3P3_MHZ_c), .D(n2659));   // src/ram.vhd(56[12:17])
    SB_DFF i5324_5325 (.Q(ram_s_221_2), .C(CLK_3P3_MHZ_c), .D(n2658));   // src/ram.vhd(56[12:17])
    SB_DFF i5321_5322 (.Q(ram_s_221_1), .C(CLK_3P3_MHZ_c), .D(n2657));   // src/ram.vhd(56[12:17])
    SB_DFF i5318_5319 (.Q(ram_s_221_0), .C(CLK_3P3_MHZ_c), .D(n2656));   // src/ram.vhd(56[12:17])
    SB_DFF i5315_5316 (.Q(ram_s_220_7), .C(CLK_3P3_MHZ_c), .D(n2655));   // src/ram.vhd(56[12:17])
    SB_DFF i5312_5313 (.Q(ram_s_220_6), .C(CLK_3P3_MHZ_c), .D(n2654));   // src/ram.vhd(56[12:17])
    SB_DFF i5309_5310 (.Q(ram_s_220_5), .C(CLK_3P3_MHZ_c), .D(n2653));   // src/ram.vhd(56[12:17])
    SB_DFF i5306_5307 (.Q(ram_s_220_4), .C(CLK_3P3_MHZ_c), .D(n2652));   // src/ram.vhd(56[12:17])
    SB_DFF i5303_5304 (.Q(ram_s_220_3), .C(CLK_3P3_MHZ_c), .D(n2651));   // src/ram.vhd(56[12:17])
    SB_DFF i5300_5301 (.Q(ram_s_220_2), .C(CLK_3P3_MHZ_c), .D(n2650));   // src/ram.vhd(56[12:17])
    SB_DFF i5297_5298 (.Q(ram_s_220_1), .C(CLK_3P3_MHZ_c), .D(n2649));   // src/ram.vhd(56[12:17])
    SB_DFF i5294_5295 (.Q(ram_s_220_0), .C(CLK_3P3_MHZ_c), .D(n2648));   // src/ram.vhd(56[12:17])
    SB_DFF i5291_5292 (.Q(ram_s_219_7), .C(CLK_3P3_MHZ_c), .D(n2647));   // src/ram.vhd(56[12:17])
    SB_DFF i5288_5289 (.Q(ram_s_219_6), .C(CLK_3P3_MHZ_c), .D(n2646));   // src/ram.vhd(56[12:17])
    SB_DFF i5285_5286 (.Q(ram_s_219_5), .C(CLK_3P3_MHZ_c), .D(n2645));   // src/ram.vhd(56[12:17])
    SB_DFF i5282_5283 (.Q(ram_s_219_4), .C(CLK_3P3_MHZ_c), .D(n2644));   // src/ram.vhd(56[12:17])
    SB_DFF i5279_5280 (.Q(ram_s_219_3), .C(CLK_3P3_MHZ_c), .D(n2643));   // src/ram.vhd(56[12:17])
    SB_DFF i5276_5277 (.Q(ram_s_219_2), .C(CLK_3P3_MHZ_c), .D(n2642));   // src/ram.vhd(56[12:17])
    SB_DFF i5273_5274 (.Q(ram_s_219_1), .C(CLK_3P3_MHZ_c), .D(n2641));   // src/ram.vhd(56[12:17])
    SB_DFF i5270_5271 (.Q(ram_s_219_0), .C(CLK_3P3_MHZ_c), .D(n2640));   // src/ram.vhd(56[12:17])
    SB_DFF i5267_5268 (.Q(ram_s_218_7), .C(CLK_3P3_MHZ_c), .D(n2639));   // src/ram.vhd(56[12:17])
    SB_DFF i5264_5265 (.Q(ram_s_218_6), .C(CLK_3P3_MHZ_c), .D(n2638));   // src/ram.vhd(56[12:17])
    SB_DFF i5261_5262 (.Q(ram_s_218_5), .C(CLK_3P3_MHZ_c), .D(n2637));   // src/ram.vhd(56[12:17])
    SB_DFF i5258_5259 (.Q(ram_s_218_4), .C(CLK_3P3_MHZ_c), .D(n2636));   // src/ram.vhd(56[12:17])
    SB_DFF i5255_5256 (.Q(ram_s_218_3), .C(CLK_3P3_MHZ_c), .D(n2635));   // src/ram.vhd(56[12:17])
    SB_DFF i5252_5253 (.Q(ram_s_218_2), .C(CLK_3P3_MHZ_c), .D(n2634));   // src/ram.vhd(56[12:17])
    SB_DFF i5249_5250 (.Q(ram_s_218_1), .C(CLK_3P3_MHZ_c), .D(n2633));   // src/ram.vhd(56[12:17])
    SB_DFF i5246_5247 (.Q(ram_s_218_0), .C(CLK_3P3_MHZ_c), .D(n2632));   // src/ram.vhd(56[12:17])
    SB_DFF i5243_5244 (.Q(ram_s_217_7), .C(CLK_3P3_MHZ_c), .D(n2631));   // src/ram.vhd(56[12:17])
    SB_DFF i5240_5241 (.Q(ram_s_217_6), .C(CLK_3P3_MHZ_c), .D(n2630));   // src/ram.vhd(56[12:17])
    SB_DFF i5237_5238 (.Q(ram_s_217_5), .C(CLK_3P3_MHZ_c), .D(n2629));   // src/ram.vhd(56[12:17])
    SB_DFF i5234_5235 (.Q(ram_s_217_4), .C(CLK_3P3_MHZ_c), .D(n2628));   // src/ram.vhd(56[12:17])
    SB_DFF i5231_5232 (.Q(ram_s_217_3), .C(CLK_3P3_MHZ_c), .D(n2627));   // src/ram.vhd(56[12:17])
    SB_DFF i5228_5229 (.Q(ram_s_217_2), .C(CLK_3P3_MHZ_c), .D(n2626));   // src/ram.vhd(56[12:17])
    SB_DFF i5225_5226 (.Q(ram_s_217_1), .C(CLK_3P3_MHZ_c), .D(n2625));   // src/ram.vhd(56[12:17])
    SB_DFF i5222_5223 (.Q(ram_s_217_0), .C(CLK_3P3_MHZ_c), .D(n2624));   // src/ram.vhd(56[12:17])
    SB_DFF i5219_5220 (.Q(ram_s_216_7), .C(CLK_3P3_MHZ_c), .D(n2623));   // src/ram.vhd(56[12:17])
    SB_DFF i5216_5217 (.Q(ram_s_216_6), .C(CLK_3P3_MHZ_c), .D(n2622));   // src/ram.vhd(56[12:17])
    SB_DFF i5213_5214 (.Q(ram_s_216_5), .C(CLK_3P3_MHZ_c), .D(n2621));   // src/ram.vhd(56[12:17])
    SB_DFF i5210_5211 (.Q(ram_s_216_4), .C(CLK_3P3_MHZ_c), .D(n2620));   // src/ram.vhd(56[12:17])
    SB_DFF i5207_5208 (.Q(ram_s_216_3), .C(CLK_3P3_MHZ_c), .D(n2619));   // src/ram.vhd(56[12:17])
    SB_DFF i5204_5205 (.Q(ram_s_216_2), .C(CLK_3P3_MHZ_c), .D(n2618));   // src/ram.vhd(56[12:17])
    SB_DFF i5201_5202 (.Q(ram_s_216_1), .C(CLK_3P3_MHZ_c), .D(n2617));   // src/ram.vhd(56[12:17])
    SB_DFF i5198_5199 (.Q(ram_s_216_0), .C(CLK_3P3_MHZ_c), .D(n2616));   // src/ram.vhd(56[12:17])
    SB_DFF i5195_5196 (.Q(ram_s_215_7), .C(CLK_3P3_MHZ_c), .D(n2615));   // src/ram.vhd(56[12:17])
    SB_DFF i5192_5193 (.Q(ram_s_215_6), .C(CLK_3P3_MHZ_c), .D(n2614));   // src/ram.vhd(56[12:17])
    SB_DFF i5189_5190 (.Q(ram_s_215_5), .C(CLK_3P3_MHZ_c), .D(n2613));   // src/ram.vhd(56[12:17])
    SB_DFF i5186_5187 (.Q(ram_s_215_4), .C(CLK_3P3_MHZ_c), .D(n2612));   // src/ram.vhd(56[12:17])
    SB_DFF i5183_5184 (.Q(ram_s_215_3), .C(CLK_3P3_MHZ_c), .D(n2611));   // src/ram.vhd(56[12:17])
    SB_DFF i5180_5181 (.Q(ram_s_215_2), .C(CLK_3P3_MHZ_c), .D(n2610));   // src/ram.vhd(56[12:17])
    SB_DFF i5177_5178 (.Q(ram_s_215_1), .C(CLK_3P3_MHZ_c), .D(n2609));   // src/ram.vhd(56[12:17])
    SB_DFF i5174_5175 (.Q(ram_s_215_0), .C(CLK_3P3_MHZ_c), .D(n2608));   // src/ram.vhd(56[12:17])
    SB_DFF i5171_5172 (.Q(ram_s_214_7), .C(CLK_3P3_MHZ_c), .D(n2607));   // src/ram.vhd(56[12:17])
    SB_DFF i5168_5169 (.Q(ram_s_214_6), .C(CLK_3P3_MHZ_c), .D(n2606));   // src/ram.vhd(56[12:17])
    SB_DFF i5165_5166 (.Q(ram_s_214_5), .C(CLK_3P3_MHZ_c), .D(n2605));   // src/ram.vhd(56[12:17])
    SB_DFF i5162_5163 (.Q(ram_s_214_4), .C(CLK_3P3_MHZ_c), .D(n2604));   // src/ram.vhd(56[12:17])
    SB_DFF i5159_5160 (.Q(ram_s_214_3), .C(CLK_3P3_MHZ_c), .D(n2603));   // src/ram.vhd(56[12:17])
    SB_DFF i5156_5157 (.Q(ram_s_214_2), .C(CLK_3P3_MHZ_c), .D(n2602));   // src/ram.vhd(56[12:17])
    SB_DFF i5153_5154 (.Q(ram_s_214_1), .C(CLK_3P3_MHZ_c), .D(n2601));   // src/ram.vhd(56[12:17])
    SB_DFF i5150_5151 (.Q(ram_s_214_0), .C(CLK_3P3_MHZ_c), .D(n2600));   // src/ram.vhd(56[12:17])
    SB_DFF i5147_5148 (.Q(ram_s_213_7), .C(CLK_3P3_MHZ_c), .D(n2599));   // src/ram.vhd(56[12:17])
    SB_DFF i5144_5145 (.Q(ram_s_213_6), .C(CLK_3P3_MHZ_c), .D(n2598));   // src/ram.vhd(56[12:17])
    SB_DFF i5141_5142 (.Q(ram_s_213_5), .C(CLK_3P3_MHZ_c), .D(n2597));   // src/ram.vhd(56[12:17])
    SB_DFF i5138_5139 (.Q(ram_s_213_4), .C(CLK_3P3_MHZ_c), .D(n2596));   // src/ram.vhd(56[12:17])
    SB_DFF i5135_5136 (.Q(ram_s_213_3), .C(CLK_3P3_MHZ_c), .D(n2595));   // src/ram.vhd(56[12:17])
    SB_DFF i5132_5133 (.Q(ram_s_213_2), .C(CLK_3P3_MHZ_c), .D(n2594));   // src/ram.vhd(56[12:17])
    SB_DFF i5129_5130 (.Q(ram_s_213_1), .C(CLK_3P3_MHZ_c), .D(n2593));   // src/ram.vhd(56[12:17])
    SB_DFF i5126_5127 (.Q(ram_s_213_0), .C(CLK_3P3_MHZ_c), .D(n2592));   // src/ram.vhd(56[12:17])
    SB_DFF i5123_5124 (.Q(ram_s_212_7), .C(CLK_3P3_MHZ_c), .D(n2591));   // src/ram.vhd(56[12:17])
    SB_DFF i5120_5121 (.Q(ram_s_212_6), .C(CLK_3P3_MHZ_c), .D(n2590));   // src/ram.vhd(56[12:17])
    SB_DFF i5117_5118 (.Q(ram_s_212_5), .C(CLK_3P3_MHZ_c), .D(n2589));   // src/ram.vhd(56[12:17])
    SB_DFF i5114_5115 (.Q(ram_s_212_4), .C(CLK_3P3_MHZ_c), .D(n2588));   // src/ram.vhd(56[12:17])
    SB_DFF i5111_5112 (.Q(ram_s_212_3), .C(CLK_3P3_MHZ_c), .D(n2587));   // src/ram.vhd(56[12:17])
    SB_DFF i5108_5109 (.Q(ram_s_212_2), .C(CLK_3P3_MHZ_c), .D(n2586));   // src/ram.vhd(56[12:17])
    SB_DFF i5105_5106 (.Q(ram_s_212_1), .C(CLK_3P3_MHZ_c), .D(n2585));   // src/ram.vhd(56[12:17])
    SB_DFF i5102_5103 (.Q(ram_s_212_0), .C(CLK_3P3_MHZ_c), .D(n2584));   // src/ram.vhd(56[12:17])
    SB_DFF i5099_5100 (.Q(ram_s_211_7), .C(CLK_3P3_MHZ_c), .D(n2583));   // src/ram.vhd(56[12:17])
    SB_DFF i5096_5097 (.Q(ram_s_211_6), .C(CLK_3P3_MHZ_c), .D(n2582));   // src/ram.vhd(56[12:17])
    SB_DFF i5093_5094 (.Q(ram_s_211_5), .C(CLK_3P3_MHZ_c), .D(n2581));   // src/ram.vhd(56[12:17])
    SB_DFF i5090_5091 (.Q(ram_s_211_4), .C(CLK_3P3_MHZ_c), .D(n2580));   // src/ram.vhd(56[12:17])
    SB_DFF i5087_5088 (.Q(ram_s_211_3), .C(CLK_3P3_MHZ_c), .D(n2579));   // src/ram.vhd(56[12:17])
    SB_DFF i5084_5085 (.Q(ram_s_211_2), .C(CLK_3P3_MHZ_c), .D(n2578));   // src/ram.vhd(56[12:17])
    SB_DFF i5081_5082 (.Q(ram_s_211_1), .C(CLK_3P3_MHZ_c), .D(n2577));   // src/ram.vhd(56[12:17])
    SB_DFF i5078_5079 (.Q(ram_s_211_0), .C(CLK_3P3_MHZ_c), .D(n2576));   // src/ram.vhd(56[12:17])
    SB_DFF i5075_5076 (.Q(ram_s_210_7), .C(CLK_3P3_MHZ_c), .D(n2575));   // src/ram.vhd(56[12:17])
    SB_DFF i5072_5073 (.Q(ram_s_210_6), .C(CLK_3P3_MHZ_c), .D(n2574));   // src/ram.vhd(56[12:17])
    SB_DFF i5069_5070 (.Q(ram_s_210_5), .C(CLK_3P3_MHZ_c), .D(n2573));   // src/ram.vhd(56[12:17])
    SB_DFF i5066_5067 (.Q(ram_s_210_4), .C(CLK_3P3_MHZ_c), .D(n2572));   // src/ram.vhd(56[12:17])
    SB_DFF i5063_5064 (.Q(ram_s_210_3), .C(CLK_3P3_MHZ_c), .D(n2571));   // src/ram.vhd(56[12:17])
    SB_DFF i5060_5061 (.Q(ram_s_210_2), .C(CLK_3P3_MHZ_c), .D(n2570));   // src/ram.vhd(56[12:17])
    SB_DFF i5057_5058 (.Q(ram_s_210_1), .C(CLK_3P3_MHZ_c), .D(n2569));   // src/ram.vhd(56[12:17])
    SB_DFF i5054_5055 (.Q(ram_s_210_0), .C(CLK_3P3_MHZ_c), .D(n2568));   // src/ram.vhd(56[12:17])
    SB_DFF i5051_5052 (.Q(ram_s_209_7), .C(CLK_3P3_MHZ_c), .D(n2567));   // src/ram.vhd(56[12:17])
    SB_DFF i5048_5049 (.Q(ram_s_209_6), .C(CLK_3P3_MHZ_c), .D(n2566));   // src/ram.vhd(56[12:17])
    SB_DFF i5045_5046 (.Q(ram_s_209_5), .C(CLK_3P3_MHZ_c), .D(n2565));   // src/ram.vhd(56[12:17])
    SB_DFF i5042_5043 (.Q(ram_s_209_4), .C(CLK_3P3_MHZ_c), .D(n2564));   // src/ram.vhd(56[12:17])
    SB_DFF i5039_5040 (.Q(ram_s_209_3), .C(CLK_3P3_MHZ_c), .D(n2563));   // src/ram.vhd(56[12:17])
    SB_DFF i5036_5037 (.Q(ram_s_209_2), .C(CLK_3P3_MHZ_c), .D(n2562));   // src/ram.vhd(56[12:17])
    SB_DFF i5033_5034 (.Q(ram_s_209_1), .C(CLK_3P3_MHZ_c), .D(n2561));   // src/ram.vhd(56[12:17])
    SB_DFF i5030_5031 (.Q(ram_s_209_0), .C(CLK_3P3_MHZ_c), .D(n2560));   // src/ram.vhd(56[12:17])
    SB_DFF i5027_5028 (.Q(ram_s_208_7), .C(CLK_3P3_MHZ_c), .D(n2559));   // src/ram.vhd(56[12:17])
    SB_DFF i5024_5025 (.Q(ram_s_208_6), .C(CLK_3P3_MHZ_c), .D(n2558));   // src/ram.vhd(56[12:17])
    SB_DFF i5021_5022 (.Q(ram_s_208_5), .C(CLK_3P3_MHZ_c), .D(n2557));   // src/ram.vhd(56[12:17])
    SB_DFF i5018_5019 (.Q(ram_s_208_4), .C(CLK_3P3_MHZ_c), .D(n2556));   // src/ram.vhd(56[12:17])
    SB_DFF i5015_5016 (.Q(ram_s_208_3), .C(CLK_3P3_MHZ_c), .D(n2555));   // src/ram.vhd(56[12:17])
    SB_DFF i5012_5013 (.Q(ram_s_208_2), .C(CLK_3P3_MHZ_c), .D(n2554));   // src/ram.vhd(56[12:17])
    SB_DFF i5009_5010 (.Q(ram_s_208_1), .C(CLK_3P3_MHZ_c), .D(n2553));   // src/ram.vhd(56[12:17])
    SB_DFF i5006_5007 (.Q(ram_s_208_0), .C(CLK_3P3_MHZ_c), .D(n2552));   // src/ram.vhd(56[12:17])
    SB_DFF i5003_5004 (.Q(ram_s_207_7), .C(CLK_3P3_MHZ_c), .D(n2551));   // src/ram.vhd(56[12:17])
    SB_DFF i5000_5001 (.Q(ram_s_207_6), .C(CLK_3P3_MHZ_c), .D(n2550));   // src/ram.vhd(56[12:17])
    SB_DFF i4997_4998 (.Q(ram_s_207_5), .C(CLK_3P3_MHZ_c), .D(n2549));   // src/ram.vhd(56[12:17])
    SB_DFF i4994_4995 (.Q(ram_s_207_4), .C(CLK_3P3_MHZ_c), .D(n2548));   // src/ram.vhd(56[12:17])
    SB_DFF i4991_4992 (.Q(ram_s_207_3), .C(CLK_3P3_MHZ_c), .D(n2547));   // src/ram.vhd(56[12:17])
    SB_DFF i4988_4989 (.Q(ram_s_207_2), .C(CLK_3P3_MHZ_c), .D(n2546));   // src/ram.vhd(56[12:17])
    SB_DFF i4985_4986 (.Q(ram_s_207_1), .C(CLK_3P3_MHZ_c), .D(n2545));   // src/ram.vhd(56[12:17])
    SB_DFF i4982_4983 (.Q(ram_s_207_0), .C(CLK_3P3_MHZ_c), .D(n2544));   // src/ram.vhd(56[12:17])
    SB_DFF i4979_4980 (.Q(ram_s_206_7), .C(CLK_3P3_MHZ_c), .D(n2543));   // src/ram.vhd(56[12:17])
    SB_DFF i4976_4977 (.Q(ram_s_206_6), .C(CLK_3P3_MHZ_c), .D(n2542));   // src/ram.vhd(56[12:17])
    SB_DFF i4973_4974 (.Q(ram_s_206_5), .C(CLK_3P3_MHZ_c), .D(n2541));   // src/ram.vhd(56[12:17])
    SB_DFF i4970_4971 (.Q(ram_s_206_4), .C(CLK_3P3_MHZ_c), .D(n2540));   // src/ram.vhd(56[12:17])
    SB_DFF i4967_4968 (.Q(ram_s_206_3), .C(CLK_3P3_MHZ_c), .D(n2539));   // src/ram.vhd(56[12:17])
    SB_DFF i4964_4965 (.Q(ram_s_206_2), .C(CLK_3P3_MHZ_c), .D(n2538));   // src/ram.vhd(56[12:17])
    SB_DFF i4961_4962 (.Q(ram_s_206_1), .C(CLK_3P3_MHZ_c), .D(n2537));   // src/ram.vhd(56[12:17])
    SB_DFF i4958_4959 (.Q(ram_s_206_0), .C(CLK_3P3_MHZ_c), .D(n2536));   // src/ram.vhd(56[12:17])
    SB_DFF i4955_4956 (.Q(ram_s_205_7), .C(CLK_3P3_MHZ_c), .D(n2535));   // src/ram.vhd(56[12:17])
    SB_DFF i4952_4953 (.Q(ram_s_205_6), .C(CLK_3P3_MHZ_c), .D(n2534));   // src/ram.vhd(56[12:17])
    SB_DFF i4949_4950 (.Q(ram_s_205_5), .C(CLK_3P3_MHZ_c), .D(n2533));   // src/ram.vhd(56[12:17])
    SB_DFF i4946_4947 (.Q(ram_s_205_4), .C(CLK_3P3_MHZ_c), .D(n2532));   // src/ram.vhd(56[12:17])
    SB_DFF i4943_4944 (.Q(ram_s_205_3), .C(CLK_3P3_MHZ_c), .D(n2531));   // src/ram.vhd(56[12:17])
    SB_DFF i4940_4941 (.Q(ram_s_205_2), .C(CLK_3P3_MHZ_c), .D(n2530));   // src/ram.vhd(56[12:17])
    SB_DFF i4937_4938 (.Q(ram_s_205_1), .C(CLK_3P3_MHZ_c), .D(n2529));   // src/ram.vhd(56[12:17])
    SB_DFF i4934_4935 (.Q(ram_s_205_0), .C(CLK_3P3_MHZ_c), .D(n2528));   // src/ram.vhd(56[12:17])
    SB_DFF i4931_4932 (.Q(ram_s_204_7), .C(CLK_3P3_MHZ_c), .D(n2527));   // src/ram.vhd(56[12:17])
    SB_DFF i4928_4929 (.Q(ram_s_204_6), .C(CLK_3P3_MHZ_c), .D(n2526));   // src/ram.vhd(56[12:17])
    SB_DFF i4925_4926 (.Q(ram_s_204_5), .C(CLK_3P3_MHZ_c), .D(n2525));   // src/ram.vhd(56[12:17])
    SB_DFF i4922_4923 (.Q(ram_s_204_4), .C(CLK_3P3_MHZ_c), .D(n2524));   // src/ram.vhd(56[12:17])
    SB_DFF i4919_4920 (.Q(ram_s_204_3), .C(CLK_3P3_MHZ_c), .D(n2523));   // src/ram.vhd(56[12:17])
    SB_DFF i4916_4917 (.Q(ram_s_204_2), .C(CLK_3P3_MHZ_c), .D(n2522));   // src/ram.vhd(56[12:17])
    SB_DFF i4913_4914 (.Q(ram_s_204_1), .C(CLK_3P3_MHZ_c), .D(n2521));   // src/ram.vhd(56[12:17])
    SB_DFF i4910_4911 (.Q(ram_s_204_0), .C(CLK_3P3_MHZ_c), .D(n2520));   // src/ram.vhd(56[12:17])
    SB_DFF i4907_4908 (.Q(ram_s_203_7), .C(CLK_3P3_MHZ_c), .D(n2519));   // src/ram.vhd(56[12:17])
    SB_DFF i4904_4905 (.Q(ram_s_203_6), .C(CLK_3P3_MHZ_c), .D(n2518));   // src/ram.vhd(56[12:17])
    SB_DFF i4901_4902 (.Q(ram_s_203_5), .C(CLK_3P3_MHZ_c), .D(n2517));   // src/ram.vhd(56[12:17])
    SB_DFF i4898_4899 (.Q(ram_s_203_4), .C(CLK_3P3_MHZ_c), .D(n2516));   // src/ram.vhd(56[12:17])
    SB_DFF i4895_4896 (.Q(ram_s_203_3), .C(CLK_3P3_MHZ_c), .D(n2515));   // src/ram.vhd(56[12:17])
    SB_DFF i4892_4893 (.Q(ram_s_203_2), .C(CLK_3P3_MHZ_c), .D(n2514));   // src/ram.vhd(56[12:17])
    SB_DFF i4889_4890 (.Q(ram_s_203_1), .C(CLK_3P3_MHZ_c), .D(n2513));   // src/ram.vhd(56[12:17])
    SB_DFF i4886_4887 (.Q(ram_s_203_0), .C(CLK_3P3_MHZ_c), .D(n2512));   // src/ram.vhd(56[12:17])
    SB_DFF i4883_4884 (.Q(ram_s_202_7), .C(CLK_3P3_MHZ_c), .D(n2511));   // src/ram.vhd(56[12:17])
    SB_DFF i4880_4881 (.Q(ram_s_202_6), .C(CLK_3P3_MHZ_c), .D(n2510));   // src/ram.vhd(56[12:17])
    SB_DFF i4877_4878 (.Q(ram_s_202_5), .C(CLK_3P3_MHZ_c), .D(n2509));   // src/ram.vhd(56[12:17])
    SB_DFF i4874_4875 (.Q(ram_s_202_4), .C(CLK_3P3_MHZ_c), .D(n2508));   // src/ram.vhd(56[12:17])
    SB_DFF i4871_4872 (.Q(ram_s_202_3), .C(CLK_3P3_MHZ_c), .D(n2507));   // src/ram.vhd(56[12:17])
    SB_DFF i4868_4869 (.Q(ram_s_202_2), .C(CLK_3P3_MHZ_c), .D(n2506));   // src/ram.vhd(56[12:17])
    SB_DFF i4865_4866 (.Q(ram_s_202_1), .C(CLK_3P3_MHZ_c), .D(n2505));   // src/ram.vhd(56[12:17])
    SB_DFF i4862_4863 (.Q(ram_s_202_0), .C(CLK_3P3_MHZ_c), .D(n2504));   // src/ram.vhd(56[12:17])
    SB_DFF i4859_4860 (.Q(ram_s_201_7), .C(CLK_3P3_MHZ_c), .D(n2503));   // src/ram.vhd(56[12:17])
    SB_DFF i4856_4857 (.Q(ram_s_201_6), .C(CLK_3P3_MHZ_c), .D(n2502));   // src/ram.vhd(56[12:17])
    SB_DFF i4853_4854 (.Q(ram_s_201_5), .C(CLK_3P3_MHZ_c), .D(n2501));   // src/ram.vhd(56[12:17])
    SB_DFF i4850_4851 (.Q(ram_s_201_4), .C(CLK_3P3_MHZ_c), .D(n2500));   // src/ram.vhd(56[12:17])
    SB_DFF i4847_4848 (.Q(ram_s_201_3), .C(CLK_3P3_MHZ_c), .D(n2499));   // src/ram.vhd(56[12:17])
    SB_DFF i4844_4845 (.Q(ram_s_201_2), .C(CLK_3P3_MHZ_c), .D(n2498));   // src/ram.vhd(56[12:17])
    SB_DFF i4841_4842 (.Q(ram_s_201_1), .C(CLK_3P3_MHZ_c), .D(n2497));   // src/ram.vhd(56[12:17])
    SB_DFF i4838_4839 (.Q(ram_s_201_0), .C(CLK_3P3_MHZ_c), .D(n2496));   // src/ram.vhd(56[12:17])
    SB_DFF i4835_4836 (.Q(ram_s_200_7), .C(CLK_3P3_MHZ_c), .D(n2495));   // src/ram.vhd(56[12:17])
    SB_DFF i4832_4833 (.Q(ram_s_200_6), .C(CLK_3P3_MHZ_c), .D(n2494));   // src/ram.vhd(56[12:17])
    SB_DFF i4829_4830 (.Q(ram_s_200_5), .C(CLK_3P3_MHZ_c), .D(n2493));   // src/ram.vhd(56[12:17])
    SB_DFF i4826_4827 (.Q(ram_s_200_4), .C(CLK_3P3_MHZ_c), .D(n2492));   // src/ram.vhd(56[12:17])
    SB_DFF i4823_4824 (.Q(ram_s_200_3), .C(CLK_3P3_MHZ_c), .D(n2491));   // src/ram.vhd(56[12:17])
    SB_DFF i4820_4821 (.Q(ram_s_200_2), .C(CLK_3P3_MHZ_c), .D(n2490));   // src/ram.vhd(56[12:17])
    SB_DFF i4817_4818 (.Q(ram_s_200_1), .C(CLK_3P3_MHZ_c), .D(n2489));   // src/ram.vhd(56[12:17])
    SB_DFF i4814_4815 (.Q(ram_s_200_0), .C(CLK_3P3_MHZ_c), .D(n2488));   // src/ram.vhd(56[12:17])
    SB_DFF i4811_4812 (.Q(ram_s_199_7), .C(CLK_3P3_MHZ_c), .D(n2487));   // src/ram.vhd(56[12:17])
    SB_DFF i4808_4809 (.Q(ram_s_199_6), .C(CLK_3P3_MHZ_c), .D(n2486));   // src/ram.vhd(56[12:17])
    SB_DFF i4805_4806 (.Q(ram_s_199_5), .C(CLK_3P3_MHZ_c), .D(n2485));   // src/ram.vhd(56[12:17])
    SB_DFF i4802_4803 (.Q(ram_s_199_4), .C(CLK_3P3_MHZ_c), .D(n2484));   // src/ram.vhd(56[12:17])
    SB_DFF i4799_4800 (.Q(ram_s_199_3), .C(CLK_3P3_MHZ_c), .D(n2483));   // src/ram.vhd(56[12:17])
    SB_DFF i4796_4797 (.Q(ram_s_199_2), .C(CLK_3P3_MHZ_c), .D(n2482));   // src/ram.vhd(56[12:17])
    SB_DFF i4793_4794 (.Q(ram_s_199_1), .C(CLK_3P3_MHZ_c), .D(n2481));   // src/ram.vhd(56[12:17])
    SB_DFF i4790_4791 (.Q(ram_s_199_0), .C(CLK_3P3_MHZ_c), .D(n2480));   // src/ram.vhd(56[12:17])
    SB_DFF i4787_4788 (.Q(ram_s_198_7), .C(CLK_3P3_MHZ_c), .D(n2479));   // src/ram.vhd(56[12:17])
    SB_DFF i4784_4785 (.Q(ram_s_198_6), .C(CLK_3P3_MHZ_c), .D(n2478));   // src/ram.vhd(56[12:17])
    SB_DFF i4781_4782 (.Q(ram_s_198_5), .C(CLK_3P3_MHZ_c), .D(n2477));   // src/ram.vhd(56[12:17])
    SB_DFF i4778_4779 (.Q(ram_s_198_4), .C(CLK_3P3_MHZ_c), .D(n2476));   // src/ram.vhd(56[12:17])
    SB_DFF i4775_4776 (.Q(ram_s_198_3), .C(CLK_3P3_MHZ_c), .D(n2475));   // src/ram.vhd(56[12:17])
    SB_DFF i4772_4773 (.Q(ram_s_198_2), .C(CLK_3P3_MHZ_c), .D(n2474));   // src/ram.vhd(56[12:17])
    SB_DFF i4769_4770 (.Q(ram_s_198_1), .C(CLK_3P3_MHZ_c), .D(n2473));   // src/ram.vhd(56[12:17])
    SB_DFF i4766_4767 (.Q(ram_s_198_0), .C(CLK_3P3_MHZ_c), .D(n2472));   // src/ram.vhd(56[12:17])
    SB_DFF i4763_4764 (.Q(ram_s_197_7), .C(CLK_3P3_MHZ_c), .D(n2471));   // src/ram.vhd(56[12:17])
    SB_DFF i4760_4761 (.Q(ram_s_197_6), .C(CLK_3P3_MHZ_c), .D(n2470));   // src/ram.vhd(56[12:17])
    SB_DFF i4757_4758 (.Q(ram_s_197_5), .C(CLK_3P3_MHZ_c), .D(n2469));   // src/ram.vhd(56[12:17])
    SB_DFF i4754_4755 (.Q(ram_s_197_4), .C(CLK_3P3_MHZ_c), .D(n2468));   // src/ram.vhd(56[12:17])
    SB_DFF i4751_4752 (.Q(ram_s_197_3), .C(CLK_3P3_MHZ_c), .D(n2467));   // src/ram.vhd(56[12:17])
    SB_DFF i4748_4749 (.Q(ram_s_197_2), .C(CLK_3P3_MHZ_c), .D(n2466));   // src/ram.vhd(56[12:17])
    SB_DFF i4745_4746 (.Q(ram_s_197_1), .C(CLK_3P3_MHZ_c), .D(n2465));   // src/ram.vhd(56[12:17])
    SB_DFF i4742_4743 (.Q(ram_s_197_0), .C(CLK_3P3_MHZ_c), .D(n2464));   // src/ram.vhd(56[12:17])
    SB_DFF i4739_4740 (.Q(ram_s_196_7), .C(CLK_3P3_MHZ_c), .D(n2463));   // src/ram.vhd(56[12:17])
    SB_DFF i4736_4737 (.Q(ram_s_196_6), .C(CLK_3P3_MHZ_c), .D(n2462));   // src/ram.vhd(56[12:17])
    SB_DFF i4733_4734 (.Q(ram_s_196_5), .C(CLK_3P3_MHZ_c), .D(n2461));   // src/ram.vhd(56[12:17])
    SB_DFF i4730_4731 (.Q(ram_s_196_4), .C(CLK_3P3_MHZ_c), .D(n2460));   // src/ram.vhd(56[12:17])
    SB_DFF i4727_4728 (.Q(ram_s_196_3), .C(CLK_3P3_MHZ_c), .D(n2459));   // src/ram.vhd(56[12:17])
    SB_DFF i4724_4725 (.Q(ram_s_196_2), .C(CLK_3P3_MHZ_c), .D(n2458));   // src/ram.vhd(56[12:17])
    SB_DFF i4721_4722 (.Q(ram_s_196_1), .C(CLK_3P3_MHZ_c), .D(n2457));   // src/ram.vhd(56[12:17])
    SB_DFF i4718_4719 (.Q(ram_s_196_0), .C(CLK_3P3_MHZ_c), .D(n2456));   // src/ram.vhd(56[12:17])
    SB_DFF i4715_4716 (.Q(ram_s_195_7), .C(CLK_3P3_MHZ_c), .D(n2455));   // src/ram.vhd(56[12:17])
    SB_DFF i4712_4713 (.Q(ram_s_195_6), .C(CLK_3P3_MHZ_c), .D(n2454));   // src/ram.vhd(56[12:17])
    SB_DFF i4709_4710 (.Q(ram_s_195_5), .C(CLK_3P3_MHZ_c), .D(n2453));   // src/ram.vhd(56[12:17])
    SB_DFF i4706_4707 (.Q(ram_s_195_4), .C(CLK_3P3_MHZ_c), .D(n2452));   // src/ram.vhd(56[12:17])
    SB_DFF i4703_4704 (.Q(ram_s_195_3), .C(CLK_3P3_MHZ_c), .D(n2451));   // src/ram.vhd(56[12:17])
    SB_DFF i4700_4701 (.Q(ram_s_195_2), .C(CLK_3P3_MHZ_c), .D(n2450));   // src/ram.vhd(56[12:17])
    SB_DFF i4697_4698 (.Q(ram_s_195_1), .C(CLK_3P3_MHZ_c), .D(n2449));   // src/ram.vhd(56[12:17])
    SB_DFF i4694_4695 (.Q(ram_s_195_0), .C(CLK_3P3_MHZ_c), .D(n2448));   // src/ram.vhd(56[12:17])
    SB_DFF i4691_4692 (.Q(ram_s_194_7), .C(CLK_3P3_MHZ_c), .D(n2447));   // src/ram.vhd(56[12:17])
    SB_DFF i4688_4689 (.Q(ram_s_194_6), .C(CLK_3P3_MHZ_c), .D(n2446));   // src/ram.vhd(56[12:17])
    SB_DFF i4685_4686 (.Q(ram_s_194_5), .C(CLK_3P3_MHZ_c), .D(n2445));   // src/ram.vhd(56[12:17])
    SB_DFF i4682_4683 (.Q(ram_s_194_4), .C(CLK_3P3_MHZ_c), .D(n2444));   // src/ram.vhd(56[12:17])
    SB_DFF i4679_4680 (.Q(ram_s_194_3), .C(CLK_3P3_MHZ_c), .D(n2443));   // src/ram.vhd(56[12:17])
    SB_DFF i4676_4677 (.Q(ram_s_194_2), .C(CLK_3P3_MHZ_c), .D(n2442));   // src/ram.vhd(56[12:17])
    SB_DFF i4673_4674 (.Q(ram_s_194_1), .C(CLK_3P3_MHZ_c), .D(n2441));   // src/ram.vhd(56[12:17])
    SB_DFF i4670_4671 (.Q(ram_s_194_0), .C(CLK_3P3_MHZ_c), .D(n2440));   // src/ram.vhd(56[12:17])
    SB_DFF i4667_4668 (.Q(ram_s_193_7), .C(CLK_3P3_MHZ_c), .D(n2439));   // src/ram.vhd(56[12:17])
    SB_DFF i4664_4665 (.Q(ram_s_193_6), .C(CLK_3P3_MHZ_c), .D(n2438));   // src/ram.vhd(56[12:17])
    SB_DFF i4661_4662 (.Q(ram_s_193_5), .C(CLK_3P3_MHZ_c), .D(n2437));   // src/ram.vhd(56[12:17])
    SB_DFF i4658_4659 (.Q(ram_s_193_4), .C(CLK_3P3_MHZ_c), .D(n2436));   // src/ram.vhd(56[12:17])
    SB_DFF i4655_4656 (.Q(ram_s_193_3), .C(CLK_3P3_MHZ_c), .D(n2435));   // src/ram.vhd(56[12:17])
    SB_DFF i4652_4653 (.Q(ram_s_193_2), .C(CLK_3P3_MHZ_c), .D(n2434));   // src/ram.vhd(56[12:17])
    SB_DFF i4649_4650 (.Q(ram_s_193_1), .C(CLK_3P3_MHZ_c), .D(n2433));   // src/ram.vhd(56[12:17])
    SB_DFF i4646_4647 (.Q(ram_s_193_0), .C(CLK_3P3_MHZ_c), .D(n2432));   // src/ram.vhd(56[12:17])
    SB_DFF i4643_4644 (.Q(ram_s_192_7), .C(CLK_3P3_MHZ_c), .D(n2431));   // src/ram.vhd(56[12:17])
    SB_DFF i4640_4641 (.Q(ram_s_192_6), .C(CLK_3P3_MHZ_c), .D(n2430));   // src/ram.vhd(56[12:17])
    SB_DFF i4637_4638 (.Q(ram_s_192_5), .C(CLK_3P3_MHZ_c), .D(n2429));   // src/ram.vhd(56[12:17])
    SB_DFF i4634_4635 (.Q(ram_s_192_4), .C(CLK_3P3_MHZ_c), .D(n2428));   // src/ram.vhd(56[12:17])
    SB_DFF i4631_4632 (.Q(ram_s_192_3), .C(CLK_3P3_MHZ_c), .D(n2427));   // src/ram.vhd(56[12:17])
    SB_DFF i4628_4629 (.Q(ram_s_192_2), .C(CLK_3P3_MHZ_c), .D(n2426));   // src/ram.vhd(56[12:17])
    SB_DFF i4625_4626 (.Q(ram_s_192_1), .C(CLK_3P3_MHZ_c), .D(n2425));   // src/ram.vhd(56[12:17])
    SB_DFF i4622_4623 (.Q(ram_s_192_0), .C(CLK_3P3_MHZ_c), .D(n2424));   // src/ram.vhd(56[12:17])
    SB_DFF i4619_4620 (.Q(ram_s_191_7), .C(CLK_3P3_MHZ_c), .D(n2423));   // src/ram.vhd(56[12:17])
    SB_DFF i4616_4617 (.Q(ram_s_191_6), .C(CLK_3P3_MHZ_c), .D(n2422));   // src/ram.vhd(56[12:17])
    SB_DFF i4613_4614 (.Q(ram_s_191_5), .C(CLK_3P3_MHZ_c), .D(n2421));   // src/ram.vhd(56[12:17])
    SB_DFF i4610_4611 (.Q(ram_s_191_4), .C(CLK_3P3_MHZ_c), .D(n2420));   // src/ram.vhd(56[12:17])
    SB_DFF i4607_4608 (.Q(ram_s_191_3), .C(CLK_3P3_MHZ_c), .D(n2419));   // src/ram.vhd(56[12:17])
    SB_DFF i4604_4605 (.Q(ram_s_191_2), .C(CLK_3P3_MHZ_c), .D(n2418));   // src/ram.vhd(56[12:17])
    SB_DFF i4601_4602 (.Q(ram_s_191_1), .C(CLK_3P3_MHZ_c), .D(n2417));   // src/ram.vhd(56[12:17])
    SB_DFF i4598_4599 (.Q(ram_s_191_0), .C(CLK_3P3_MHZ_c), .D(n2416));   // src/ram.vhd(56[12:17])
    SB_DFF i4595_4596 (.Q(ram_s_190_7), .C(CLK_3P3_MHZ_c), .D(n2415));   // src/ram.vhd(56[12:17])
    SB_DFF i4592_4593 (.Q(ram_s_190_6), .C(CLK_3P3_MHZ_c), .D(n2414));   // src/ram.vhd(56[12:17])
    SB_DFF i4589_4590 (.Q(ram_s_190_5), .C(CLK_3P3_MHZ_c), .D(n2413));   // src/ram.vhd(56[12:17])
    SB_DFF i4586_4587 (.Q(ram_s_190_4), .C(CLK_3P3_MHZ_c), .D(n2412));   // src/ram.vhd(56[12:17])
    SB_DFF i4583_4584 (.Q(ram_s_190_3), .C(CLK_3P3_MHZ_c), .D(n2411));   // src/ram.vhd(56[12:17])
    SB_DFF i4580_4581 (.Q(ram_s_190_2), .C(CLK_3P3_MHZ_c), .D(n2410));   // src/ram.vhd(56[12:17])
    SB_DFF i4577_4578 (.Q(ram_s_190_1), .C(CLK_3P3_MHZ_c), .D(n2409));   // src/ram.vhd(56[12:17])
    SB_DFF i4574_4575 (.Q(ram_s_190_0), .C(CLK_3P3_MHZ_c), .D(n2408));   // src/ram.vhd(56[12:17])
    SB_DFF i4571_4572 (.Q(ram_s_189_7), .C(CLK_3P3_MHZ_c), .D(n2407));   // src/ram.vhd(56[12:17])
    SB_DFF i4568_4569 (.Q(ram_s_189_6), .C(CLK_3P3_MHZ_c), .D(n2406));   // src/ram.vhd(56[12:17])
    SB_DFF i4565_4566 (.Q(ram_s_189_5), .C(CLK_3P3_MHZ_c), .D(n2405));   // src/ram.vhd(56[12:17])
    SB_DFF i4562_4563 (.Q(ram_s_189_4), .C(CLK_3P3_MHZ_c), .D(n2404));   // src/ram.vhd(56[12:17])
    SB_DFF i4559_4560 (.Q(ram_s_189_3), .C(CLK_3P3_MHZ_c), .D(n2403));   // src/ram.vhd(56[12:17])
    SB_DFF i4556_4557 (.Q(ram_s_189_2), .C(CLK_3P3_MHZ_c), .D(n2402));   // src/ram.vhd(56[12:17])
    SB_DFF i4553_4554 (.Q(ram_s_189_1), .C(CLK_3P3_MHZ_c), .D(n2401));   // src/ram.vhd(56[12:17])
    SB_DFF i4550_4551 (.Q(ram_s_189_0), .C(CLK_3P3_MHZ_c), .D(n2400));   // src/ram.vhd(56[12:17])
    SB_DFF i4547_4548 (.Q(ram_s_188_7), .C(CLK_3P3_MHZ_c), .D(n2399));   // src/ram.vhd(56[12:17])
    SB_DFF i4544_4545 (.Q(ram_s_188_6), .C(CLK_3P3_MHZ_c), .D(n2398));   // src/ram.vhd(56[12:17])
    SB_DFF i4541_4542 (.Q(ram_s_188_5), .C(CLK_3P3_MHZ_c), .D(n2397));   // src/ram.vhd(56[12:17])
    SB_DFF i4538_4539 (.Q(ram_s_188_4), .C(CLK_3P3_MHZ_c), .D(n2396));   // src/ram.vhd(56[12:17])
    SB_DFF i4535_4536 (.Q(ram_s_188_3), .C(CLK_3P3_MHZ_c), .D(n2395));   // src/ram.vhd(56[12:17])
    SB_DFF i4532_4533 (.Q(ram_s_188_2), .C(CLK_3P3_MHZ_c), .D(n2394));   // src/ram.vhd(56[12:17])
    SB_DFF i4529_4530 (.Q(ram_s_188_1), .C(CLK_3P3_MHZ_c), .D(n2393));   // src/ram.vhd(56[12:17])
    SB_DFF i4526_4527 (.Q(ram_s_188_0), .C(CLK_3P3_MHZ_c), .D(n2392));   // src/ram.vhd(56[12:17])
    SB_DFF i4523_4524 (.Q(ram_s_187_7), .C(CLK_3P3_MHZ_c), .D(n2391));   // src/ram.vhd(56[12:17])
    SB_DFF i4520_4521 (.Q(ram_s_187_6), .C(CLK_3P3_MHZ_c), .D(n2390));   // src/ram.vhd(56[12:17])
    SB_DFF i4517_4518 (.Q(ram_s_187_5), .C(CLK_3P3_MHZ_c), .D(n2389));   // src/ram.vhd(56[12:17])
    SB_DFF i4514_4515 (.Q(ram_s_187_4), .C(CLK_3P3_MHZ_c), .D(n2388));   // src/ram.vhd(56[12:17])
    SB_DFF i4511_4512 (.Q(ram_s_187_3), .C(CLK_3P3_MHZ_c), .D(n2387));   // src/ram.vhd(56[12:17])
    SB_DFF i4508_4509 (.Q(ram_s_187_2), .C(CLK_3P3_MHZ_c), .D(n2386));   // src/ram.vhd(56[12:17])
    SB_DFF i4505_4506 (.Q(ram_s_187_1), .C(CLK_3P3_MHZ_c), .D(n2385));   // src/ram.vhd(56[12:17])
    SB_DFF i4502_4503 (.Q(ram_s_187_0), .C(CLK_3P3_MHZ_c), .D(n2384));   // src/ram.vhd(56[12:17])
    SB_DFF i4499_4500 (.Q(ram_s_186_7), .C(CLK_3P3_MHZ_c), .D(n2383));   // src/ram.vhd(56[12:17])
    SB_DFF i4496_4497 (.Q(ram_s_186_6), .C(CLK_3P3_MHZ_c), .D(n2382));   // src/ram.vhd(56[12:17])
    SB_DFF i4493_4494 (.Q(ram_s_186_5), .C(CLK_3P3_MHZ_c), .D(n2381));   // src/ram.vhd(56[12:17])
    SB_DFF i4490_4491 (.Q(ram_s_186_4), .C(CLK_3P3_MHZ_c), .D(n2380));   // src/ram.vhd(56[12:17])
    SB_DFF i4487_4488 (.Q(ram_s_186_3), .C(CLK_3P3_MHZ_c), .D(n2379));   // src/ram.vhd(56[12:17])
    SB_DFF i4484_4485 (.Q(ram_s_186_2), .C(CLK_3P3_MHZ_c), .D(n2378));   // src/ram.vhd(56[12:17])
    SB_DFF i4481_4482 (.Q(ram_s_186_1), .C(CLK_3P3_MHZ_c), .D(n2377));   // src/ram.vhd(56[12:17])
    SB_DFF i4478_4479 (.Q(ram_s_186_0), .C(CLK_3P3_MHZ_c), .D(n2376));   // src/ram.vhd(56[12:17])
    SB_DFF i4475_4476 (.Q(ram_s_185_7), .C(CLK_3P3_MHZ_c), .D(n2375));   // src/ram.vhd(56[12:17])
    SB_DFF i4472_4473 (.Q(ram_s_185_6), .C(CLK_3P3_MHZ_c), .D(n2374));   // src/ram.vhd(56[12:17])
    SB_DFF i4469_4470 (.Q(ram_s_185_5), .C(CLK_3P3_MHZ_c), .D(n2373));   // src/ram.vhd(56[12:17])
    SB_DFF i4466_4467 (.Q(ram_s_185_4), .C(CLK_3P3_MHZ_c), .D(n2372));   // src/ram.vhd(56[12:17])
    SB_DFF i4463_4464 (.Q(ram_s_185_3), .C(CLK_3P3_MHZ_c), .D(n2371));   // src/ram.vhd(56[12:17])
    SB_DFF i4460_4461 (.Q(ram_s_185_2), .C(CLK_3P3_MHZ_c), .D(n2370));   // src/ram.vhd(56[12:17])
    SB_DFF i4457_4458 (.Q(ram_s_185_1), .C(CLK_3P3_MHZ_c), .D(n2369));   // src/ram.vhd(56[12:17])
    SB_DFF i4454_4455 (.Q(ram_s_185_0), .C(CLK_3P3_MHZ_c), .D(n2368));   // src/ram.vhd(56[12:17])
    SB_DFF i4451_4452 (.Q(ram_s_184_7), .C(CLK_3P3_MHZ_c), .D(n2367));   // src/ram.vhd(56[12:17])
    SB_DFF i4448_4449 (.Q(ram_s_184_6), .C(CLK_3P3_MHZ_c), .D(n2366));   // src/ram.vhd(56[12:17])
    SB_DFF i4445_4446 (.Q(ram_s_184_5), .C(CLK_3P3_MHZ_c), .D(n2365));   // src/ram.vhd(56[12:17])
    SB_DFF i4442_4443 (.Q(ram_s_184_4), .C(CLK_3P3_MHZ_c), .D(n2364));   // src/ram.vhd(56[12:17])
    SB_DFF i4439_4440 (.Q(ram_s_184_3), .C(CLK_3P3_MHZ_c), .D(n2363));   // src/ram.vhd(56[12:17])
    SB_DFF i4436_4437 (.Q(ram_s_184_2), .C(CLK_3P3_MHZ_c), .D(n2362));   // src/ram.vhd(56[12:17])
    SB_DFF i4433_4434 (.Q(ram_s_184_1), .C(CLK_3P3_MHZ_c), .D(n2361));   // src/ram.vhd(56[12:17])
    SB_DFF i4430_4431 (.Q(ram_s_184_0), .C(CLK_3P3_MHZ_c), .D(n2360));   // src/ram.vhd(56[12:17])
    SB_DFF i4427_4428 (.Q(ram_s_183_7), .C(CLK_3P3_MHZ_c), .D(n2359));   // src/ram.vhd(56[12:17])
    SB_DFF i4424_4425 (.Q(ram_s_183_6), .C(CLK_3P3_MHZ_c), .D(n2358));   // src/ram.vhd(56[12:17])
    SB_DFF i4421_4422 (.Q(ram_s_183_5), .C(CLK_3P3_MHZ_c), .D(n2357));   // src/ram.vhd(56[12:17])
    SB_DFF i4418_4419 (.Q(ram_s_183_4), .C(CLK_3P3_MHZ_c), .D(n2356));   // src/ram.vhd(56[12:17])
    SB_DFF i4415_4416 (.Q(ram_s_183_3), .C(CLK_3P3_MHZ_c), .D(n2355));   // src/ram.vhd(56[12:17])
    SB_DFF i4412_4413 (.Q(ram_s_183_2), .C(CLK_3P3_MHZ_c), .D(n2354));   // src/ram.vhd(56[12:17])
    SB_DFF i4409_4410 (.Q(ram_s_183_1), .C(CLK_3P3_MHZ_c), .D(n2353));   // src/ram.vhd(56[12:17])
    SB_DFF i4406_4407 (.Q(ram_s_183_0), .C(CLK_3P3_MHZ_c), .D(n2352));   // src/ram.vhd(56[12:17])
    SB_DFF i4403_4404 (.Q(ram_s_182_7), .C(CLK_3P3_MHZ_c), .D(n2351));   // src/ram.vhd(56[12:17])
    SB_DFF i4400_4401 (.Q(ram_s_182_6), .C(CLK_3P3_MHZ_c), .D(n2350));   // src/ram.vhd(56[12:17])
    SB_DFF i4397_4398 (.Q(ram_s_182_5), .C(CLK_3P3_MHZ_c), .D(n2349));   // src/ram.vhd(56[12:17])
    SB_DFF i4394_4395 (.Q(ram_s_182_4), .C(CLK_3P3_MHZ_c), .D(n2348));   // src/ram.vhd(56[12:17])
    SB_DFF i4391_4392 (.Q(ram_s_182_3), .C(CLK_3P3_MHZ_c), .D(n2347));   // src/ram.vhd(56[12:17])
    SB_DFF i4388_4389 (.Q(ram_s_182_2), .C(CLK_3P3_MHZ_c), .D(n2346));   // src/ram.vhd(56[12:17])
    SB_DFF i4385_4386 (.Q(ram_s_182_1), .C(CLK_3P3_MHZ_c), .D(n2345));   // src/ram.vhd(56[12:17])
    SB_DFF i4382_4383 (.Q(ram_s_182_0), .C(CLK_3P3_MHZ_c), .D(n2344));   // src/ram.vhd(56[12:17])
    SB_DFF i4379_4380 (.Q(ram_s_181_7), .C(CLK_3P3_MHZ_c), .D(n2343));   // src/ram.vhd(56[12:17])
    SB_DFF i4376_4377 (.Q(ram_s_181_6), .C(CLK_3P3_MHZ_c), .D(n2342));   // src/ram.vhd(56[12:17])
    SB_DFF i4373_4374 (.Q(ram_s_181_5), .C(CLK_3P3_MHZ_c), .D(n2341));   // src/ram.vhd(56[12:17])
    SB_DFF i4370_4371 (.Q(ram_s_181_4), .C(CLK_3P3_MHZ_c), .D(n2340));   // src/ram.vhd(56[12:17])
    SB_DFF i4367_4368 (.Q(ram_s_181_3), .C(CLK_3P3_MHZ_c), .D(n2339));   // src/ram.vhd(56[12:17])
    SB_DFF i4364_4365 (.Q(ram_s_181_2), .C(CLK_3P3_MHZ_c), .D(n2338));   // src/ram.vhd(56[12:17])
    SB_DFF i4361_4362 (.Q(ram_s_181_1), .C(CLK_3P3_MHZ_c), .D(n2337));   // src/ram.vhd(56[12:17])
    SB_DFF i4358_4359 (.Q(ram_s_181_0), .C(CLK_3P3_MHZ_c), .D(n2336));   // src/ram.vhd(56[12:17])
    SB_DFF i4355_4356 (.Q(ram_s_180_7), .C(CLK_3P3_MHZ_c), .D(n2335));   // src/ram.vhd(56[12:17])
    SB_DFF i4352_4353 (.Q(ram_s_180_6), .C(CLK_3P3_MHZ_c), .D(n2334));   // src/ram.vhd(56[12:17])
    SB_DFF i4349_4350 (.Q(ram_s_180_5), .C(CLK_3P3_MHZ_c), .D(n2333));   // src/ram.vhd(56[12:17])
    SB_DFF i4346_4347 (.Q(ram_s_180_4), .C(CLK_3P3_MHZ_c), .D(n2332));   // src/ram.vhd(56[12:17])
    SB_DFF i4343_4344 (.Q(ram_s_180_3), .C(CLK_3P3_MHZ_c), .D(n2331));   // src/ram.vhd(56[12:17])
    SB_DFF i4340_4341 (.Q(ram_s_180_2), .C(CLK_3P3_MHZ_c), .D(n2330));   // src/ram.vhd(56[12:17])
    SB_DFF i4337_4338 (.Q(ram_s_180_1), .C(CLK_3P3_MHZ_c), .D(n2329));   // src/ram.vhd(56[12:17])
    SB_DFF i4334_4335 (.Q(ram_s_180_0), .C(CLK_3P3_MHZ_c), .D(n2328));   // src/ram.vhd(56[12:17])
    SB_DFF i4331_4332 (.Q(ram_s_179_7), .C(CLK_3P3_MHZ_c), .D(n2327));   // src/ram.vhd(56[12:17])
    SB_DFF i4328_4329 (.Q(ram_s_179_6), .C(CLK_3P3_MHZ_c), .D(n2326));   // src/ram.vhd(56[12:17])
    SB_DFF i4325_4326 (.Q(ram_s_179_5), .C(CLK_3P3_MHZ_c), .D(n2325));   // src/ram.vhd(56[12:17])
    SB_DFF i4322_4323 (.Q(ram_s_179_4), .C(CLK_3P3_MHZ_c), .D(n2324));   // src/ram.vhd(56[12:17])
    SB_DFF i4319_4320 (.Q(ram_s_179_3), .C(CLK_3P3_MHZ_c), .D(n2323));   // src/ram.vhd(56[12:17])
    SB_DFF i4316_4317 (.Q(ram_s_179_2), .C(CLK_3P3_MHZ_c), .D(n2322));   // src/ram.vhd(56[12:17])
    SB_DFF i4313_4314 (.Q(ram_s_179_1), .C(CLK_3P3_MHZ_c), .D(n2321));   // src/ram.vhd(56[12:17])
    SB_DFF i4310_4311 (.Q(ram_s_179_0), .C(CLK_3P3_MHZ_c), .D(n2320));   // src/ram.vhd(56[12:17])
    SB_DFF i4307_4308 (.Q(ram_s_178_7), .C(CLK_3P3_MHZ_c), .D(n2319));   // src/ram.vhd(56[12:17])
    SB_DFF i4304_4305 (.Q(ram_s_178_6), .C(CLK_3P3_MHZ_c), .D(n2318));   // src/ram.vhd(56[12:17])
    SB_DFF i4301_4302 (.Q(ram_s_178_5), .C(CLK_3P3_MHZ_c), .D(n2317));   // src/ram.vhd(56[12:17])
    SB_DFF i4298_4299 (.Q(ram_s_178_4), .C(CLK_3P3_MHZ_c), .D(n2316));   // src/ram.vhd(56[12:17])
    SB_DFF i4295_4296 (.Q(ram_s_178_3), .C(CLK_3P3_MHZ_c), .D(n2315));   // src/ram.vhd(56[12:17])
    SB_DFF i4292_4293 (.Q(ram_s_178_2), .C(CLK_3P3_MHZ_c), .D(n2314));   // src/ram.vhd(56[12:17])
    SB_DFF i4289_4290 (.Q(ram_s_178_1), .C(CLK_3P3_MHZ_c), .D(n2313));   // src/ram.vhd(56[12:17])
    SB_DFF i4286_4287 (.Q(ram_s_178_0), .C(CLK_3P3_MHZ_c), .D(n2312));   // src/ram.vhd(56[12:17])
    SB_DFF i4283_4284 (.Q(ram_s_177_7), .C(CLK_3P3_MHZ_c), .D(n2311));   // src/ram.vhd(56[12:17])
    SB_DFF i4280_4281 (.Q(ram_s_177_6), .C(CLK_3P3_MHZ_c), .D(n2310));   // src/ram.vhd(56[12:17])
    SB_DFF i4277_4278 (.Q(ram_s_177_5), .C(CLK_3P3_MHZ_c), .D(n2309));   // src/ram.vhd(56[12:17])
    SB_DFF i4274_4275 (.Q(ram_s_177_4), .C(CLK_3P3_MHZ_c), .D(n2308));   // src/ram.vhd(56[12:17])
    SB_DFF i4271_4272 (.Q(ram_s_177_3), .C(CLK_3P3_MHZ_c), .D(n2307));   // src/ram.vhd(56[12:17])
    SB_DFF i4268_4269 (.Q(ram_s_177_2), .C(CLK_3P3_MHZ_c), .D(n2306));   // src/ram.vhd(56[12:17])
    SB_DFF i4265_4266 (.Q(ram_s_177_1), .C(CLK_3P3_MHZ_c), .D(n2305));   // src/ram.vhd(56[12:17])
    SB_DFF i4262_4263 (.Q(ram_s_177_0), .C(CLK_3P3_MHZ_c), .D(n2304));   // src/ram.vhd(56[12:17])
    SB_DFF i4259_4260 (.Q(ram_s_176_7), .C(CLK_3P3_MHZ_c), .D(n2303));   // src/ram.vhd(56[12:17])
    SB_DFF i4256_4257 (.Q(ram_s_176_6), .C(CLK_3P3_MHZ_c), .D(n2302));   // src/ram.vhd(56[12:17])
    SB_DFF i4253_4254 (.Q(ram_s_176_5), .C(CLK_3P3_MHZ_c), .D(n2301));   // src/ram.vhd(56[12:17])
    SB_DFF i4250_4251 (.Q(ram_s_176_4), .C(CLK_3P3_MHZ_c), .D(n2300));   // src/ram.vhd(56[12:17])
    SB_DFF i4247_4248 (.Q(ram_s_176_3), .C(CLK_3P3_MHZ_c), .D(n2299));   // src/ram.vhd(56[12:17])
    SB_DFF i4244_4245 (.Q(ram_s_176_2), .C(CLK_3P3_MHZ_c), .D(n2298));   // src/ram.vhd(56[12:17])
    SB_DFF i4241_4242 (.Q(ram_s_176_1), .C(CLK_3P3_MHZ_c), .D(n2297));   // src/ram.vhd(56[12:17])
    SB_DFF i4238_4239 (.Q(ram_s_176_0), .C(CLK_3P3_MHZ_c), .D(n2296));   // src/ram.vhd(56[12:17])
    SB_DFF i4235_4236 (.Q(ram_s_175_7), .C(CLK_3P3_MHZ_c), .D(n2295));   // src/ram.vhd(56[12:17])
    SB_DFF i4232_4233 (.Q(ram_s_175_6), .C(CLK_3P3_MHZ_c), .D(n2294));   // src/ram.vhd(56[12:17])
    SB_DFF i4229_4230 (.Q(ram_s_175_5), .C(CLK_3P3_MHZ_c), .D(n2293));   // src/ram.vhd(56[12:17])
    SB_DFF i4226_4227 (.Q(ram_s_175_4), .C(CLK_3P3_MHZ_c), .D(n2292));   // src/ram.vhd(56[12:17])
    SB_DFF i4223_4224 (.Q(ram_s_175_3), .C(CLK_3P3_MHZ_c), .D(n2291));   // src/ram.vhd(56[12:17])
    SB_DFF i4220_4221 (.Q(ram_s_175_2), .C(CLK_3P3_MHZ_c), .D(n2290));   // src/ram.vhd(56[12:17])
    SB_DFF i4217_4218 (.Q(ram_s_175_1), .C(CLK_3P3_MHZ_c), .D(n2289));   // src/ram.vhd(56[12:17])
    SB_DFF i4214_4215 (.Q(ram_s_175_0), .C(CLK_3P3_MHZ_c), .D(n2288));   // src/ram.vhd(56[12:17])
    SB_DFF i4211_4212 (.Q(ram_s_174_7), .C(CLK_3P3_MHZ_c), .D(n2287));   // src/ram.vhd(56[12:17])
    SB_DFF i4208_4209 (.Q(ram_s_174_6), .C(CLK_3P3_MHZ_c), .D(n2286));   // src/ram.vhd(56[12:17])
    SB_DFF i4205_4206 (.Q(ram_s_174_5), .C(CLK_3P3_MHZ_c), .D(n2285));   // src/ram.vhd(56[12:17])
    SB_DFF i4202_4203 (.Q(ram_s_174_4), .C(CLK_3P3_MHZ_c), .D(n2284));   // src/ram.vhd(56[12:17])
    SB_DFF i4199_4200 (.Q(ram_s_174_3), .C(CLK_3P3_MHZ_c), .D(n2283));   // src/ram.vhd(56[12:17])
    SB_DFF i4196_4197 (.Q(ram_s_174_2), .C(CLK_3P3_MHZ_c), .D(n2282));   // src/ram.vhd(56[12:17])
    SB_DFF i4193_4194 (.Q(ram_s_174_1), .C(CLK_3P3_MHZ_c), .D(n2281));   // src/ram.vhd(56[12:17])
    SB_DFF i4190_4191 (.Q(ram_s_174_0), .C(CLK_3P3_MHZ_c), .D(n2280));   // src/ram.vhd(56[12:17])
    SB_DFF i4187_4188 (.Q(ram_s_173_7), .C(CLK_3P3_MHZ_c), .D(n2279));   // src/ram.vhd(56[12:17])
    SB_DFF i4184_4185 (.Q(ram_s_173_6), .C(CLK_3P3_MHZ_c), .D(n2278));   // src/ram.vhd(56[12:17])
    SB_DFF i4181_4182 (.Q(ram_s_173_5), .C(CLK_3P3_MHZ_c), .D(n2277));   // src/ram.vhd(56[12:17])
    SB_DFF i4178_4179 (.Q(ram_s_173_4), .C(CLK_3P3_MHZ_c), .D(n2276));   // src/ram.vhd(56[12:17])
    SB_DFF i4175_4176 (.Q(ram_s_173_3), .C(CLK_3P3_MHZ_c), .D(n2275));   // src/ram.vhd(56[12:17])
    SB_DFF i4172_4173 (.Q(ram_s_173_2), .C(CLK_3P3_MHZ_c), .D(n2274));   // src/ram.vhd(56[12:17])
    SB_DFF i4169_4170 (.Q(ram_s_173_1), .C(CLK_3P3_MHZ_c), .D(n2273));   // src/ram.vhd(56[12:17])
    SB_DFF i4166_4167 (.Q(ram_s_173_0), .C(CLK_3P3_MHZ_c), .D(n2272));   // src/ram.vhd(56[12:17])
    SB_DFF i4163_4164 (.Q(ram_s_172_7), .C(CLK_3P3_MHZ_c), .D(n2271));   // src/ram.vhd(56[12:17])
    SB_DFF i4160_4161 (.Q(ram_s_172_6), .C(CLK_3P3_MHZ_c), .D(n2270));   // src/ram.vhd(56[12:17])
    SB_DFF i4157_4158 (.Q(ram_s_172_5), .C(CLK_3P3_MHZ_c), .D(n2269));   // src/ram.vhd(56[12:17])
    SB_DFF i4154_4155 (.Q(ram_s_172_4), .C(CLK_3P3_MHZ_c), .D(n2268));   // src/ram.vhd(56[12:17])
    SB_DFF i4151_4152 (.Q(ram_s_172_3), .C(CLK_3P3_MHZ_c), .D(n2267));   // src/ram.vhd(56[12:17])
    SB_DFF i4148_4149 (.Q(ram_s_172_2), .C(CLK_3P3_MHZ_c), .D(n2266));   // src/ram.vhd(56[12:17])
    SB_DFF i4145_4146 (.Q(ram_s_172_1), .C(CLK_3P3_MHZ_c), .D(n2265));   // src/ram.vhd(56[12:17])
    SB_DFF i4142_4143 (.Q(ram_s_172_0), .C(CLK_3P3_MHZ_c), .D(n2264));   // src/ram.vhd(56[12:17])
    SB_DFF i4139_4140 (.Q(ram_s_171_7), .C(CLK_3P3_MHZ_c), .D(n2263));   // src/ram.vhd(56[12:17])
    SB_DFF i4136_4137 (.Q(ram_s_171_6), .C(CLK_3P3_MHZ_c), .D(n2262));   // src/ram.vhd(56[12:17])
    SB_DFF i4133_4134 (.Q(ram_s_171_5), .C(CLK_3P3_MHZ_c), .D(n2261));   // src/ram.vhd(56[12:17])
    SB_DFF i4130_4131 (.Q(ram_s_171_4), .C(CLK_3P3_MHZ_c), .D(n2260));   // src/ram.vhd(56[12:17])
    SB_DFF i4127_4128 (.Q(ram_s_171_3), .C(CLK_3P3_MHZ_c), .D(n2259));   // src/ram.vhd(56[12:17])
    SB_DFF i4124_4125 (.Q(ram_s_171_2), .C(CLK_3P3_MHZ_c), .D(n2258));   // src/ram.vhd(56[12:17])
    SB_DFF i4121_4122 (.Q(ram_s_171_1), .C(CLK_3P3_MHZ_c), .D(n2257));   // src/ram.vhd(56[12:17])
    SB_DFF i4118_4119 (.Q(ram_s_171_0), .C(CLK_3P3_MHZ_c), .D(n2256));   // src/ram.vhd(56[12:17])
    SB_DFF i4115_4116 (.Q(ram_s_170_7), .C(CLK_3P3_MHZ_c), .D(n2255));   // src/ram.vhd(56[12:17])
    SB_DFF i4112_4113 (.Q(ram_s_170_6), .C(CLK_3P3_MHZ_c), .D(n2254));   // src/ram.vhd(56[12:17])
    SB_DFF i4109_4110 (.Q(ram_s_170_5), .C(CLK_3P3_MHZ_c), .D(n2253));   // src/ram.vhd(56[12:17])
    SB_DFF i4106_4107 (.Q(ram_s_170_4), .C(CLK_3P3_MHZ_c), .D(n2252));   // src/ram.vhd(56[12:17])
    SB_DFF i4103_4104 (.Q(ram_s_170_3), .C(CLK_3P3_MHZ_c), .D(n2251));   // src/ram.vhd(56[12:17])
    SB_DFF i4100_4101 (.Q(ram_s_170_2), .C(CLK_3P3_MHZ_c), .D(n2250));   // src/ram.vhd(56[12:17])
    SB_DFF i4097_4098 (.Q(ram_s_170_1), .C(CLK_3P3_MHZ_c), .D(n2249));   // src/ram.vhd(56[12:17])
    SB_DFF i4094_4095 (.Q(ram_s_170_0), .C(CLK_3P3_MHZ_c), .D(n2248));   // src/ram.vhd(56[12:17])
    SB_DFF i4091_4092 (.Q(ram_s_169_7), .C(CLK_3P3_MHZ_c), .D(n2247));   // src/ram.vhd(56[12:17])
    SB_DFF i4088_4089 (.Q(ram_s_169_6), .C(CLK_3P3_MHZ_c), .D(n2246));   // src/ram.vhd(56[12:17])
    SB_DFF i4085_4086 (.Q(ram_s_169_5), .C(CLK_3P3_MHZ_c), .D(n2245));   // src/ram.vhd(56[12:17])
    SB_DFF i4082_4083 (.Q(ram_s_169_4), .C(CLK_3P3_MHZ_c), .D(n2244));   // src/ram.vhd(56[12:17])
    SB_DFF i4079_4080 (.Q(ram_s_169_3), .C(CLK_3P3_MHZ_c), .D(n2243));   // src/ram.vhd(56[12:17])
    SB_DFF i4076_4077 (.Q(ram_s_169_2), .C(CLK_3P3_MHZ_c), .D(n2242));   // src/ram.vhd(56[12:17])
    SB_DFF i4073_4074 (.Q(ram_s_169_1), .C(CLK_3P3_MHZ_c), .D(n2241));   // src/ram.vhd(56[12:17])
    SB_DFF i4070_4071 (.Q(ram_s_169_0), .C(CLK_3P3_MHZ_c), .D(n2240));   // src/ram.vhd(56[12:17])
    SB_DFF i4067_4068 (.Q(ram_s_168_7), .C(CLK_3P3_MHZ_c), .D(n2239));   // src/ram.vhd(56[12:17])
    SB_DFF i4064_4065 (.Q(ram_s_168_6), .C(CLK_3P3_MHZ_c), .D(n2238));   // src/ram.vhd(56[12:17])
    SB_DFF i4061_4062 (.Q(ram_s_168_5), .C(CLK_3P3_MHZ_c), .D(n2237));   // src/ram.vhd(56[12:17])
    SB_DFF i4058_4059 (.Q(ram_s_168_4), .C(CLK_3P3_MHZ_c), .D(n2236));   // src/ram.vhd(56[12:17])
    SB_DFF i4055_4056 (.Q(ram_s_168_3), .C(CLK_3P3_MHZ_c), .D(n2235));   // src/ram.vhd(56[12:17])
    SB_DFF i4052_4053 (.Q(ram_s_168_2), .C(CLK_3P3_MHZ_c), .D(n2234));   // src/ram.vhd(56[12:17])
    SB_DFF i4049_4050 (.Q(ram_s_168_1), .C(CLK_3P3_MHZ_c), .D(n2233));   // src/ram.vhd(56[12:17])
    SB_DFF i4046_4047 (.Q(ram_s_168_0), .C(CLK_3P3_MHZ_c), .D(n2232));   // src/ram.vhd(56[12:17])
    SB_DFF i4043_4044 (.Q(ram_s_167_7), .C(CLK_3P3_MHZ_c), .D(n2231));   // src/ram.vhd(56[12:17])
    SB_DFF i4040_4041 (.Q(ram_s_167_6), .C(CLK_3P3_MHZ_c), .D(n2230));   // src/ram.vhd(56[12:17])
    SB_DFF i4037_4038 (.Q(ram_s_167_5), .C(CLK_3P3_MHZ_c), .D(n2229));   // src/ram.vhd(56[12:17])
    SB_DFF i4034_4035 (.Q(ram_s_167_4), .C(CLK_3P3_MHZ_c), .D(n2228));   // src/ram.vhd(56[12:17])
    SB_DFF i4031_4032 (.Q(ram_s_167_3), .C(CLK_3P3_MHZ_c), .D(n2227));   // src/ram.vhd(56[12:17])
    SB_DFF i4028_4029 (.Q(ram_s_167_2), .C(CLK_3P3_MHZ_c), .D(n2226));   // src/ram.vhd(56[12:17])
    SB_DFF i4025_4026 (.Q(ram_s_167_1), .C(CLK_3P3_MHZ_c), .D(n2225));   // src/ram.vhd(56[12:17])
    SB_DFF i4022_4023 (.Q(ram_s_167_0), .C(CLK_3P3_MHZ_c), .D(n2224));   // src/ram.vhd(56[12:17])
    SB_DFF i4019_4020 (.Q(ram_s_166_7), .C(CLK_3P3_MHZ_c), .D(n2223));   // src/ram.vhd(56[12:17])
    SB_DFF i4016_4017 (.Q(ram_s_166_6), .C(CLK_3P3_MHZ_c), .D(n2222));   // src/ram.vhd(56[12:17])
    SB_DFF i4013_4014 (.Q(ram_s_166_5), .C(CLK_3P3_MHZ_c), .D(n2221));   // src/ram.vhd(56[12:17])
    SB_DFF i4010_4011 (.Q(ram_s_166_4), .C(CLK_3P3_MHZ_c), .D(n2220));   // src/ram.vhd(56[12:17])
    SB_DFF i4007_4008 (.Q(ram_s_166_3), .C(CLK_3P3_MHZ_c), .D(n2219));   // src/ram.vhd(56[12:17])
    SB_DFF i4004_4005 (.Q(ram_s_166_2), .C(CLK_3P3_MHZ_c), .D(n2218));   // src/ram.vhd(56[12:17])
    SB_DFF i4001_4002 (.Q(ram_s_166_1), .C(CLK_3P3_MHZ_c), .D(n2217));   // src/ram.vhd(56[12:17])
    SB_DFF i3998_3999 (.Q(ram_s_166_0), .C(CLK_3P3_MHZ_c), .D(n2216));   // src/ram.vhd(56[12:17])
    SB_DFF i3995_3996 (.Q(ram_s_165_7), .C(CLK_3P3_MHZ_c), .D(n2215));   // src/ram.vhd(56[12:17])
    SB_DFF i3992_3993 (.Q(ram_s_165_6), .C(CLK_3P3_MHZ_c), .D(n2214));   // src/ram.vhd(56[12:17])
    SB_DFF i3989_3990 (.Q(ram_s_165_5), .C(CLK_3P3_MHZ_c), .D(n2213));   // src/ram.vhd(56[12:17])
    SB_DFF i3986_3987 (.Q(ram_s_165_4), .C(CLK_3P3_MHZ_c), .D(n2212));   // src/ram.vhd(56[12:17])
    SB_DFF i3983_3984 (.Q(ram_s_165_3), .C(CLK_3P3_MHZ_c), .D(n2211));   // src/ram.vhd(56[12:17])
    SB_DFF i3980_3981 (.Q(ram_s_165_2), .C(CLK_3P3_MHZ_c), .D(n2210));   // src/ram.vhd(56[12:17])
    SB_DFF i3977_3978 (.Q(ram_s_165_1), .C(CLK_3P3_MHZ_c), .D(n2209));   // src/ram.vhd(56[12:17])
    SB_DFF i3974_3975 (.Q(ram_s_165_0), .C(CLK_3P3_MHZ_c), .D(n2208));   // src/ram.vhd(56[12:17])
    SB_DFF i3971_3972 (.Q(ram_s_164_7), .C(CLK_3P3_MHZ_c), .D(n2207));   // src/ram.vhd(56[12:17])
    SB_DFF i3968_3969 (.Q(ram_s_164_6), .C(CLK_3P3_MHZ_c), .D(n2206));   // src/ram.vhd(56[12:17])
    SB_DFF i3965_3966 (.Q(ram_s_164_5), .C(CLK_3P3_MHZ_c), .D(n2205));   // src/ram.vhd(56[12:17])
    SB_DFF i3962_3963 (.Q(ram_s_164_4), .C(CLK_3P3_MHZ_c), .D(n2204));   // src/ram.vhd(56[12:17])
    SB_DFF i3959_3960 (.Q(ram_s_164_3), .C(CLK_3P3_MHZ_c), .D(n2203));   // src/ram.vhd(56[12:17])
    SB_DFF i3956_3957 (.Q(ram_s_164_2), .C(CLK_3P3_MHZ_c), .D(n2202));   // src/ram.vhd(56[12:17])
    SB_DFF i3953_3954 (.Q(ram_s_164_1), .C(CLK_3P3_MHZ_c), .D(n2201));   // src/ram.vhd(56[12:17])
    SB_DFF i3950_3951 (.Q(ram_s_164_0), .C(CLK_3P3_MHZ_c), .D(n2200));   // src/ram.vhd(56[12:17])
    SB_DFF i3947_3948 (.Q(ram_s_163_7), .C(CLK_3P3_MHZ_c), .D(n2199));   // src/ram.vhd(56[12:17])
    SB_DFF i3944_3945 (.Q(ram_s_163_6), .C(CLK_3P3_MHZ_c), .D(n2198));   // src/ram.vhd(56[12:17])
    SB_DFF i3941_3942 (.Q(ram_s_163_5), .C(CLK_3P3_MHZ_c), .D(n2197));   // src/ram.vhd(56[12:17])
    SB_DFF i3938_3939 (.Q(ram_s_163_4), .C(CLK_3P3_MHZ_c), .D(n2196));   // src/ram.vhd(56[12:17])
    SB_DFF i3935_3936 (.Q(ram_s_163_3), .C(CLK_3P3_MHZ_c), .D(n2195));   // src/ram.vhd(56[12:17])
    SB_DFF i3932_3933 (.Q(ram_s_163_2), .C(CLK_3P3_MHZ_c), .D(n2194));   // src/ram.vhd(56[12:17])
    SB_DFF i3929_3930 (.Q(ram_s_163_1), .C(CLK_3P3_MHZ_c), .D(n2193));   // src/ram.vhd(56[12:17])
    SB_DFF i3926_3927 (.Q(ram_s_163_0), .C(CLK_3P3_MHZ_c), .D(n2192));   // src/ram.vhd(56[12:17])
    SB_DFF i3923_3924 (.Q(ram_s_162_7), .C(CLK_3P3_MHZ_c), .D(n2191));   // src/ram.vhd(56[12:17])
    SB_DFF i3920_3921 (.Q(ram_s_162_6), .C(CLK_3P3_MHZ_c), .D(n2190));   // src/ram.vhd(56[12:17])
    SB_DFF i3917_3918 (.Q(ram_s_162_5), .C(CLK_3P3_MHZ_c), .D(n2189));   // src/ram.vhd(56[12:17])
    SB_DFF i3914_3915 (.Q(ram_s_162_4), .C(CLK_3P3_MHZ_c), .D(n2188));   // src/ram.vhd(56[12:17])
    SB_DFF i3911_3912 (.Q(ram_s_162_3), .C(CLK_3P3_MHZ_c), .D(n2187));   // src/ram.vhd(56[12:17])
    SB_DFF i3908_3909 (.Q(ram_s_162_2), .C(CLK_3P3_MHZ_c), .D(n2186));   // src/ram.vhd(56[12:17])
    SB_DFF i3905_3906 (.Q(ram_s_162_1), .C(CLK_3P3_MHZ_c), .D(n2185));   // src/ram.vhd(56[12:17])
    SB_DFF i3902_3903 (.Q(ram_s_162_0), .C(CLK_3P3_MHZ_c), .D(n2184));   // src/ram.vhd(56[12:17])
    SB_DFF i3899_3900 (.Q(ram_s_161_7), .C(CLK_3P3_MHZ_c), .D(n2183));   // src/ram.vhd(56[12:17])
    SB_DFF i3896_3897 (.Q(ram_s_161_6), .C(CLK_3P3_MHZ_c), .D(n2182));   // src/ram.vhd(56[12:17])
    SB_DFF i3893_3894 (.Q(ram_s_161_5), .C(CLK_3P3_MHZ_c), .D(n2181));   // src/ram.vhd(56[12:17])
    SB_DFF i3890_3891 (.Q(ram_s_161_4), .C(CLK_3P3_MHZ_c), .D(n2180));   // src/ram.vhd(56[12:17])
    SB_DFF i3887_3888 (.Q(ram_s_161_3), .C(CLK_3P3_MHZ_c), .D(n2179));   // src/ram.vhd(56[12:17])
    SB_DFF i3884_3885 (.Q(ram_s_161_2), .C(CLK_3P3_MHZ_c), .D(n2178));   // src/ram.vhd(56[12:17])
    SB_DFF i3881_3882 (.Q(ram_s_161_1), .C(CLK_3P3_MHZ_c), .D(n2177));   // src/ram.vhd(56[12:17])
    SB_DFF i3878_3879 (.Q(ram_s_161_0), .C(CLK_3P3_MHZ_c), .D(n2176));   // src/ram.vhd(56[12:17])
    SB_DFF i3875_3876 (.Q(ram_s_160_7), .C(CLK_3P3_MHZ_c), .D(n2175));   // src/ram.vhd(56[12:17])
    SB_DFF i3872_3873 (.Q(ram_s_160_6), .C(CLK_3P3_MHZ_c), .D(n2174));   // src/ram.vhd(56[12:17])
    SB_DFF i3869_3870 (.Q(ram_s_160_5), .C(CLK_3P3_MHZ_c), .D(n2173));   // src/ram.vhd(56[12:17])
    SB_DFF i3866_3867 (.Q(ram_s_160_4), .C(CLK_3P3_MHZ_c), .D(n2172));   // src/ram.vhd(56[12:17])
    SB_DFF i3863_3864 (.Q(ram_s_160_3), .C(CLK_3P3_MHZ_c), .D(n2171));   // src/ram.vhd(56[12:17])
    SB_DFF i3860_3861 (.Q(ram_s_160_2), .C(CLK_3P3_MHZ_c), .D(n2170));   // src/ram.vhd(56[12:17])
    SB_DFF i3857_3858 (.Q(ram_s_160_1), .C(CLK_3P3_MHZ_c), .D(n2169));   // src/ram.vhd(56[12:17])
    SB_DFF i3854_3855 (.Q(ram_s_160_0), .C(CLK_3P3_MHZ_c), .D(n2168));   // src/ram.vhd(56[12:17])
    SB_DFF i3851_3852 (.Q(ram_s_159_7), .C(CLK_3P3_MHZ_c), .D(n2167));   // src/ram.vhd(56[12:17])
    SB_DFF i3848_3849 (.Q(ram_s_159_6), .C(CLK_3P3_MHZ_c), .D(n2166));   // src/ram.vhd(56[12:17])
    SB_DFF i3845_3846 (.Q(ram_s_159_5), .C(CLK_3P3_MHZ_c), .D(n2165));   // src/ram.vhd(56[12:17])
    SB_DFF i3842_3843 (.Q(ram_s_159_4), .C(CLK_3P3_MHZ_c), .D(n2164));   // src/ram.vhd(56[12:17])
    SB_DFF i3839_3840 (.Q(ram_s_159_3), .C(CLK_3P3_MHZ_c), .D(n2163));   // src/ram.vhd(56[12:17])
    SB_DFF i3836_3837 (.Q(ram_s_159_2), .C(CLK_3P3_MHZ_c), .D(n2162));   // src/ram.vhd(56[12:17])
    SB_DFF i3833_3834 (.Q(ram_s_159_1), .C(CLK_3P3_MHZ_c), .D(n2161));   // src/ram.vhd(56[12:17])
    SB_DFF i3830_3831 (.Q(ram_s_159_0), .C(CLK_3P3_MHZ_c), .D(n2160));   // src/ram.vhd(56[12:17])
    SB_DFF i3827_3828 (.Q(ram_s_158_7), .C(CLK_3P3_MHZ_c), .D(n2159));   // src/ram.vhd(56[12:17])
    SB_DFF i3824_3825 (.Q(ram_s_158_6), .C(CLK_3P3_MHZ_c), .D(n2158));   // src/ram.vhd(56[12:17])
    SB_DFF i3821_3822 (.Q(ram_s_158_5), .C(CLK_3P3_MHZ_c), .D(n2157));   // src/ram.vhd(56[12:17])
    SB_DFF i3818_3819 (.Q(ram_s_158_4), .C(CLK_3P3_MHZ_c), .D(n2156));   // src/ram.vhd(56[12:17])
    SB_DFF i3815_3816 (.Q(ram_s_158_3), .C(CLK_3P3_MHZ_c), .D(n2155));   // src/ram.vhd(56[12:17])
    SB_DFF i3812_3813 (.Q(ram_s_158_2), .C(CLK_3P3_MHZ_c), .D(n2154));   // src/ram.vhd(56[12:17])
    SB_DFF i3809_3810 (.Q(ram_s_158_1), .C(CLK_3P3_MHZ_c), .D(n2153));   // src/ram.vhd(56[12:17])
    SB_DFF i3806_3807 (.Q(ram_s_158_0), .C(CLK_3P3_MHZ_c), .D(n2152));   // src/ram.vhd(56[12:17])
    SB_DFF i3803_3804 (.Q(ram_s_157_7), .C(CLK_3P3_MHZ_c), .D(n2151));   // src/ram.vhd(56[12:17])
    SB_DFF i3800_3801 (.Q(ram_s_157_6), .C(CLK_3P3_MHZ_c), .D(n2150));   // src/ram.vhd(56[12:17])
    SB_DFF i3797_3798 (.Q(ram_s_157_5), .C(CLK_3P3_MHZ_c), .D(n2149));   // src/ram.vhd(56[12:17])
    SB_DFF i3794_3795 (.Q(ram_s_157_4), .C(CLK_3P3_MHZ_c), .D(n2148));   // src/ram.vhd(56[12:17])
    SB_DFF i3791_3792 (.Q(ram_s_157_3), .C(CLK_3P3_MHZ_c), .D(n2147));   // src/ram.vhd(56[12:17])
    SB_DFF i3788_3789 (.Q(ram_s_157_2), .C(CLK_3P3_MHZ_c), .D(n2146));   // src/ram.vhd(56[12:17])
    SB_DFF i3785_3786 (.Q(ram_s_157_1), .C(CLK_3P3_MHZ_c), .D(n2145));   // src/ram.vhd(56[12:17])
    SB_DFF i3782_3783 (.Q(ram_s_157_0), .C(CLK_3P3_MHZ_c), .D(n2144));   // src/ram.vhd(56[12:17])
    SB_DFF i3779_3780 (.Q(ram_s_156_7), .C(CLK_3P3_MHZ_c), .D(n2143));   // src/ram.vhd(56[12:17])
    SB_DFF i3776_3777 (.Q(ram_s_156_6), .C(CLK_3P3_MHZ_c), .D(n2142));   // src/ram.vhd(56[12:17])
    SB_DFF i3773_3774 (.Q(ram_s_156_5), .C(CLK_3P3_MHZ_c), .D(n2141));   // src/ram.vhd(56[12:17])
    SB_DFF i3770_3771 (.Q(ram_s_156_4), .C(CLK_3P3_MHZ_c), .D(n2140));   // src/ram.vhd(56[12:17])
    SB_DFF i3767_3768 (.Q(ram_s_156_3), .C(CLK_3P3_MHZ_c), .D(n2139));   // src/ram.vhd(56[12:17])
    SB_DFF i3764_3765 (.Q(ram_s_156_2), .C(CLK_3P3_MHZ_c), .D(n2138));   // src/ram.vhd(56[12:17])
    SB_DFF i3761_3762 (.Q(ram_s_156_1), .C(CLK_3P3_MHZ_c), .D(n2137));   // src/ram.vhd(56[12:17])
    SB_DFF i3758_3759 (.Q(ram_s_156_0), .C(CLK_3P3_MHZ_c), .D(n2136));   // src/ram.vhd(56[12:17])
    SB_DFF i3755_3756 (.Q(ram_s_155_7), .C(CLK_3P3_MHZ_c), .D(n2135));   // src/ram.vhd(56[12:17])
    SB_DFF i3752_3753 (.Q(ram_s_155_6), .C(CLK_3P3_MHZ_c), .D(n2134));   // src/ram.vhd(56[12:17])
    SB_DFF i3749_3750 (.Q(ram_s_155_5), .C(CLK_3P3_MHZ_c), .D(n2133));   // src/ram.vhd(56[12:17])
    SB_DFF i3746_3747 (.Q(ram_s_155_4), .C(CLK_3P3_MHZ_c), .D(n2132));   // src/ram.vhd(56[12:17])
    SB_DFF i3743_3744 (.Q(ram_s_155_3), .C(CLK_3P3_MHZ_c), .D(n2131));   // src/ram.vhd(56[12:17])
    SB_DFF i3740_3741 (.Q(ram_s_155_2), .C(CLK_3P3_MHZ_c), .D(n2130));   // src/ram.vhd(56[12:17])
    SB_DFF i3737_3738 (.Q(ram_s_155_1), .C(CLK_3P3_MHZ_c), .D(n2129));   // src/ram.vhd(56[12:17])
    SB_DFF i3734_3735 (.Q(ram_s_155_0), .C(CLK_3P3_MHZ_c), .D(n2128));   // src/ram.vhd(56[12:17])
    SB_DFF i3731_3732 (.Q(ram_s_154_7), .C(CLK_3P3_MHZ_c), .D(n2127));   // src/ram.vhd(56[12:17])
    SB_DFF i3728_3729 (.Q(ram_s_154_6), .C(CLK_3P3_MHZ_c), .D(n2126));   // src/ram.vhd(56[12:17])
    SB_DFF i3725_3726 (.Q(ram_s_154_5), .C(CLK_3P3_MHZ_c), .D(n2125));   // src/ram.vhd(56[12:17])
    SB_DFF i3722_3723 (.Q(ram_s_154_4), .C(CLK_3P3_MHZ_c), .D(n2124));   // src/ram.vhd(56[12:17])
    SB_DFF i3719_3720 (.Q(ram_s_154_3), .C(CLK_3P3_MHZ_c), .D(n2123));   // src/ram.vhd(56[12:17])
    SB_DFF i3716_3717 (.Q(ram_s_154_2), .C(CLK_3P3_MHZ_c), .D(n2122));   // src/ram.vhd(56[12:17])
    SB_DFF i3713_3714 (.Q(ram_s_154_1), .C(CLK_3P3_MHZ_c), .D(n2121));   // src/ram.vhd(56[12:17])
    SB_DFF i3710_3711 (.Q(ram_s_154_0), .C(CLK_3P3_MHZ_c), .D(n2120));   // src/ram.vhd(56[12:17])
    SB_DFF i3707_3708 (.Q(ram_s_153_7), .C(CLK_3P3_MHZ_c), .D(n2119));   // src/ram.vhd(56[12:17])
    SB_DFF i3704_3705 (.Q(ram_s_153_6), .C(CLK_3P3_MHZ_c), .D(n2118));   // src/ram.vhd(56[12:17])
    SB_DFF i3701_3702 (.Q(ram_s_153_5), .C(CLK_3P3_MHZ_c), .D(n2117));   // src/ram.vhd(56[12:17])
    SB_DFF i3698_3699 (.Q(ram_s_153_4), .C(CLK_3P3_MHZ_c), .D(n2116));   // src/ram.vhd(56[12:17])
    SB_DFF i3695_3696 (.Q(ram_s_153_3), .C(CLK_3P3_MHZ_c), .D(n2115));   // src/ram.vhd(56[12:17])
    SB_DFF i3692_3693 (.Q(ram_s_153_2), .C(CLK_3P3_MHZ_c), .D(n2114));   // src/ram.vhd(56[12:17])
    SB_DFF i3689_3690 (.Q(ram_s_153_1), .C(CLK_3P3_MHZ_c), .D(n2113));   // src/ram.vhd(56[12:17])
    SB_DFF i3686_3687 (.Q(ram_s_153_0), .C(CLK_3P3_MHZ_c), .D(n2112));   // src/ram.vhd(56[12:17])
    SB_DFF i3683_3684 (.Q(ram_s_152_7), .C(CLK_3P3_MHZ_c), .D(n2111));   // src/ram.vhd(56[12:17])
    SB_DFF i3680_3681 (.Q(ram_s_152_6), .C(CLK_3P3_MHZ_c), .D(n2110));   // src/ram.vhd(56[12:17])
    SB_DFF i3677_3678 (.Q(ram_s_152_5), .C(CLK_3P3_MHZ_c), .D(n2109));   // src/ram.vhd(56[12:17])
    SB_DFF i3674_3675 (.Q(ram_s_152_4), .C(CLK_3P3_MHZ_c), .D(n2108));   // src/ram.vhd(56[12:17])
    SB_DFF i3671_3672 (.Q(ram_s_152_3), .C(CLK_3P3_MHZ_c), .D(n2107));   // src/ram.vhd(56[12:17])
    SB_DFF i3668_3669 (.Q(ram_s_152_2), .C(CLK_3P3_MHZ_c), .D(n2106));   // src/ram.vhd(56[12:17])
    SB_DFF i3665_3666 (.Q(ram_s_152_1), .C(CLK_3P3_MHZ_c), .D(n2105));   // src/ram.vhd(56[12:17])
    SB_DFF i3662_3663 (.Q(ram_s_152_0), .C(CLK_3P3_MHZ_c), .D(n2104));   // src/ram.vhd(56[12:17])
    SB_DFF i3659_3660 (.Q(ram_s_151_7), .C(CLK_3P3_MHZ_c), .D(n2103));   // src/ram.vhd(56[12:17])
    SB_DFF i3656_3657 (.Q(ram_s_151_6), .C(CLK_3P3_MHZ_c), .D(n2102));   // src/ram.vhd(56[12:17])
    SB_DFF i3653_3654 (.Q(ram_s_151_5), .C(CLK_3P3_MHZ_c), .D(n2101));   // src/ram.vhd(56[12:17])
    SB_DFF i3650_3651 (.Q(ram_s_151_4), .C(CLK_3P3_MHZ_c), .D(n2100));   // src/ram.vhd(56[12:17])
    SB_DFF i3647_3648 (.Q(ram_s_151_3), .C(CLK_3P3_MHZ_c), .D(n2099));   // src/ram.vhd(56[12:17])
    SB_DFF i3644_3645 (.Q(ram_s_151_2), .C(CLK_3P3_MHZ_c), .D(n2098));   // src/ram.vhd(56[12:17])
    SB_DFF i3641_3642 (.Q(ram_s_151_1), .C(CLK_3P3_MHZ_c), .D(n2097));   // src/ram.vhd(56[12:17])
    SB_DFF i3638_3639 (.Q(ram_s_151_0), .C(CLK_3P3_MHZ_c), .D(n2096));   // src/ram.vhd(56[12:17])
    SB_DFF i3635_3636 (.Q(ram_s_150_7), .C(CLK_3P3_MHZ_c), .D(n2095));   // src/ram.vhd(56[12:17])
    SB_DFF i3632_3633 (.Q(ram_s_150_6), .C(CLK_3P3_MHZ_c), .D(n2094));   // src/ram.vhd(56[12:17])
    SB_DFF i3629_3630 (.Q(ram_s_150_5), .C(CLK_3P3_MHZ_c), .D(n2093));   // src/ram.vhd(56[12:17])
    SB_DFF i3626_3627 (.Q(ram_s_150_4), .C(CLK_3P3_MHZ_c), .D(n2092));   // src/ram.vhd(56[12:17])
    SB_DFF i3623_3624 (.Q(ram_s_150_3), .C(CLK_3P3_MHZ_c), .D(n2091));   // src/ram.vhd(56[12:17])
    SB_DFF i3620_3621 (.Q(ram_s_150_2), .C(CLK_3P3_MHZ_c), .D(n2090));   // src/ram.vhd(56[12:17])
    SB_DFF i3617_3618 (.Q(ram_s_150_1), .C(CLK_3P3_MHZ_c), .D(n2089));   // src/ram.vhd(56[12:17])
    SB_DFF i3614_3615 (.Q(ram_s_150_0), .C(CLK_3P3_MHZ_c), .D(n2088));   // src/ram.vhd(56[12:17])
    SB_DFF i3611_3612 (.Q(ram_s_149_7), .C(CLK_3P3_MHZ_c), .D(n2087));   // src/ram.vhd(56[12:17])
    SB_DFF i3608_3609 (.Q(ram_s_149_6), .C(CLK_3P3_MHZ_c), .D(n2086));   // src/ram.vhd(56[12:17])
    SB_DFF i3605_3606 (.Q(ram_s_149_5), .C(CLK_3P3_MHZ_c), .D(n2085));   // src/ram.vhd(56[12:17])
    SB_DFF i3602_3603 (.Q(ram_s_149_4), .C(CLK_3P3_MHZ_c), .D(n2084));   // src/ram.vhd(56[12:17])
    SB_DFF i3599_3600 (.Q(ram_s_149_3), .C(CLK_3P3_MHZ_c), .D(n2083));   // src/ram.vhd(56[12:17])
    SB_DFF i3596_3597 (.Q(ram_s_149_2), .C(CLK_3P3_MHZ_c), .D(n2082));   // src/ram.vhd(56[12:17])
    SB_DFF i3593_3594 (.Q(ram_s_149_1), .C(CLK_3P3_MHZ_c), .D(n2081));   // src/ram.vhd(56[12:17])
    SB_DFF i3590_3591 (.Q(ram_s_149_0), .C(CLK_3P3_MHZ_c), .D(n2080));   // src/ram.vhd(56[12:17])
    SB_DFF i3587_3588 (.Q(ram_s_148_7), .C(CLK_3P3_MHZ_c), .D(n2079));   // src/ram.vhd(56[12:17])
    SB_DFF i3584_3585 (.Q(ram_s_148_6), .C(CLK_3P3_MHZ_c), .D(n2078));   // src/ram.vhd(56[12:17])
    SB_DFF i3581_3582 (.Q(ram_s_148_5), .C(CLK_3P3_MHZ_c), .D(n2077));   // src/ram.vhd(56[12:17])
    SB_DFF i3578_3579 (.Q(ram_s_148_4), .C(CLK_3P3_MHZ_c), .D(n2076));   // src/ram.vhd(56[12:17])
    SB_DFF i3575_3576 (.Q(ram_s_148_3), .C(CLK_3P3_MHZ_c), .D(n2075));   // src/ram.vhd(56[12:17])
    SB_DFF i3572_3573 (.Q(ram_s_148_2), .C(CLK_3P3_MHZ_c), .D(n2074));   // src/ram.vhd(56[12:17])
    SB_DFF i3569_3570 (.Q(ram_s_148_1), .C(CLK_3P3_MHZ_c), .D(n2073));   // src/ram.vhd(56[12:17])
    SB_DFF i3566_3567 (.Q(ram_s_148_0), .C(CLK_3P3_MHZ_c), .D(n2072));   // src/ram.vhd(56[12:17])
    SB_DFF i3563_3564 (.Q(ram_s_147_7), .C(CLK_3P3_MHZ_c), .D(n2071));   // src/ram.vhd(56[12:17])
    SB_DFF i3560_3561 (.Q(ram_s_147_6), .C(CLK_3P3_MHZ_c), .D(n2070));   // src/ram.vhd(56[12:17])
    SB_DFF i3557_3558 (.Q(ram_s_147_5), .C(CLK_3P3_MHZ_c), .D(n2069));   // src/ram.vhd(56[12:17])
    SB_DFF i3554_3555 (.Q(ram_s_147_4), .C(CLK_3P3_MHZ_c), .D(n2068));   // src/ram.vhd(56[12:17])
    SB_DFF i3551_3552 (.Q(ram_s_147_3), .C(CLK_3P3_MHZ_c), .D(n2067));   // src/ram.vhd(56[12:17])
    SB_DFF i3548_3549 (.Q(ram_s_147_2), .C(CLK_3P3_MHZ_c), .D(n2066));   // src/ram.vhd(56[12:17])
    SB_DFF i3545_3546 (.Q(ram_s_147_1), .C(CLK_3P3_MHZ_c), .D(n2065));   // src/ram.vhd(56[12:17])
    SB_DFF i3542_3543 (.Q(ram_s_147_0), .C(CLK_3P3_MHZ_c), .D(n2064));   // src/ram.vhd(56[12:17])
    SB_DFF i3539_3540 (.Q(ram_s_146_7), .C(CLK_3P3_MHZ_c), .D(n2063));   // src/ram.vhd(56[12:17])
    SB_DFF i3536_3537 (.Q(ram_s_146_6), .C(CLK_3P3_MHZ_c), .D(n2062));   // src/ram.vhd(56[12:17])
    SB_DFF i3533_3534 (.Q(ram_s_146_5), .C(CLK_3P3_MHZ_c), .D(n2061));   // src/ram.vhd(56[12:17])
    SB_DFF i3530_3531 (.Q(ram_s_146_4), .C(CLK_3P3_MHZ_c), .D(n2060));   // src/ram.vhd(56[12:17])
    SB_DFF i3527_3528 (.Q(ram_s_146_3), .C(CLK_3P3_MHZ_c), .D(n2059));   // src/ram.vhd(56[12:17])
    SB_DFF i3524_3525 (.Q(ram_s_146_2), .C(CLK_3P3_MHZ_c), .D(n2058));   // src/ram.vhd(56[12:17])
    SB_DFF i3521_3522 (.Q(ram_s_146_1), .C(CLK_3P3_MHZ_c), .D(n2057));   // src/ram.vhd(56[12:17])
    SB_DFF i3518_3519 (.Q(ram_s_146_0), .C(CLK_3P3_MHZ_c), .D(n2056));   // src/ram.vhd(56[12:17])
    SB_DFF i3515_3516 (.Q(ram_s_145_7), .C(CLK_3P3_MHZ_c), .D(n2055));   // src/ram.vhd(56[12:17])
    SB_DFF i3512_3513 (.Q(ram_s_145_6), .C(CLK_3P3_MHZ_c), .D(n2054));   // src/ram.vhd(56[12:17])
    SB_DFF i3509_3510 (.Q(ram_s_145_5), .C(CLK_3P3_MHZ_c), .D(n2053));   // src/ram.vhd(56[12:17])
    SB_DFF i3506_3507 (.Q(ram_s_145_4), .C(CLK_3P3_MHZ_c), .D(n2052));   // src/ram.vhd(56[12:17])
    SB_DFF i3503_3504 (.Q(ram_s_145_3), .C(CLK_3P3_MHZ_c), .D(n2051));   // src/ram.vhd(56[12:17])
    SB_DFF i3500_3501 (.Q(ram_s_145_2), .C(CLK_3P3_MHZ_c), .D(n2050));   // src/ram.vhd(56[12:17])
    SB_DFF i3497_3498 (.Q(ram_s_145_1), .C(CLK_3P3_MHZ_c), .D(n2049));   // src/ram.vhd(56[12:17])
    SB_DFF i3494_3495 (.Q(ram_s_145_0), .C(CLK_3P3_MHZ_c), .D(n2048));   // src/ram.vhd(56[12:17])
    SB_DFF i3491_3492 (.Q(ram_s_144_7), .C(CLK_3P3_MHZ_c), .D(n2047));   // src/ram.vhd(56[12:17])
    SB_DFF i3488_3489 (.Q(ram_s_144_6), .C(CLK_3P3_MHZ_c), .D(n2046));   // src/ram.vhd(56[12:17])
    SB_DFF i3485_3486 (.Q(ram_s_144_5), .C(CLK_3P3_MHZ_c), .D(n2045));   // src/ram.vhd(56[12:17])
    SB_DFF i3482_3483 (.Q(ram_s_144_4), .C(CLK_3P3_MHZ_c), .D(n2044));   // src/ram.vhd(56[12:17])
    SB_DFF i3479_3480 (.Q(ram_s_144_3), .C(CLK_3P3_MHZ_c), .D(n2043));   // src/ram.vhd(56[12:17])
    SB_DFF i3476_3477 (.Q(ram_s_144_2), .C(CLK_3P3_MHZ_c), .D(n2042));   // src/ram.vhd(56[12:17])
    SB_DFF i3473_3474 (.Q(ram_s_144_1), .C(CLK_3P3_MHZ_c), .D(n2041));   // src/ram.vhd(56[12:17])
    SB_DFF i3470_3471 (.Q(ram_s_144_0), .C(CLK_3P3_MHZ_c), .D(n2040));   // src/ram.vhd(56[12:17])
    SB_DFF i3467_3468 (.Q(ram_s_143_7), .C(CLK_3P3_MHZ_c), .D(n2039));   // src/ram.vhd(56[12:17])
    SB_DFF i3464_3465 (.Q(ram_s_143_6), .C(CLK_3P3_MHZ_c), .D(n2038));   // src/ram.vhd(56[12:17])
    SB_DFF i3461_3462 (.Q(ram_s_143_5), .C(CLK_3P3_MHZ_c), .D(n2037));   // src/ram.vhd(56[12:17])
    SB_DFF i3458_3459 (.Q(ram_s_143_4), .C(CLK_3P3_MHZ_c), .D(n2036));   // src/ram.vhd(56[12:17])
    SB_DFF i3455_3456 (.Q(ram_s_143_3), .C(CLK_3P3_MHZ_c), .D(n2035));   // src/ram.vhd(56[12:17])
    SB_DFF i3452_3453 (.Q(ram_s_143_2), .C(CLK_3P3_MHZ_c), .D(n2034));   // src/ram.vhd(56[12:17])
    SB_DFF i3449_3450 (.Q(ram_s_143_1), .C(CLK_3P3_MHZ_c), .D(n2033));   // src/ram.vhd(56[12:17])
    SB_DFF i3446_3447 (.Q(ram_s_143_0), .C(CLK_3P3_MHZ_c), .D(n2032));   // src/ram.vhd(56[12:17])
    SB_DFF i3443_3444 (.Q(ram_s_142_7), .C(CLK_3P3_MHZ_c), .D(n2031));   // src/ram.vhd(56[12:17])
    SB_DFF i3440_3441 (.Q(ram_s_142_6), .C(CLK_3P3_MHZ_c), .D(n2030));   // src/ram.vhd(56[12:17])
    SB_DFF i3437_3438 (.Q(ram_s_142_5), .C(CLK_3P3_MHZ_c), .D(n2029));   // src/ram.vhd(56[12:17])
    SB_DFF i3434_3435 (.Q(ram_s_142_4), .C(CLK_3P3_MHZ_c), .D(n2028));   // src/ram.vhd(56[12:17])
    SB_DFF i3431_3432 (.Q(ram_s_142_3), .C(CLK_3P3_MHZ_c), .D(n2027));   // src/ram.vhd(56[12:17])
    SB_DFF i3428_3429 (.Q(ram_s_142_2), .C(CLK_3P3_MHZ_c), .D(n2026));   // src/ram.vhd(56[12:17])
    SB_DFF i3425_3426 (.Q(ram_s_142_1), .C(CLK_3P3_MHZ_c), .D(n2025));   // src/ram.vhd(56[12:17])
    SB_DFF i3422_3423 (.Q(ram_s_142_0), .C(CLK_3P3_MHZ_c), .D(n2024));   // src/ram.vhd(56[12:17])
    SB_DFF i3419_3420 (.Q(ram_s_141_7), .C(CLK_3P3_MHZ_c), .D(n2023));   // src/ram.vhd(56[12:17])
    SB_DFF i3416_3417 (.Q(ram_s_141_6), .C(CLK_3P3_MHZ_c), .D(n2022));   // src/ram.vhd(56[12:17])
    SB_DFF i3413_3414 (.Q(ram_s_141_5), .C(CLK_3P3_MHZ_c), .D(n2021));   // src/ram.vhd(56[12:17])
    SB_DFF i3410_3411 (.Q(ram_s_141_4), .C(CLK_3P3_MHZ_c), .D(n2020));   // src/ram.vhd(56[12:17])
    SB_DFF i3407_3408 (.Q(ram_s_141_3), .C(CLK_3P3_MHZ_c), .D(n2019));   // src/ram.vhd(56[12:17])
    SB_DFF i3404_3405 (.Q(ram_s_141_2), .C(CLK_3P3_MHZ_c), .D(n2018));   // src/ram.vhd(56[12:17])
    SB_DFF i3401_3402 (.Q(ram_s_141_1), .C(CLK_3P3_MHZ_c), .D(n2017));   // src/ram.vhd(56[12:17])
    SB_DFF i3398_3399 (.Q(ram_s_141_0), .C(CLK_3P3_MHZ_c), .D(n2016));   // src/ram.vhd(56[12:17])
    SB_DFF i3395_3396 (.Q(ram_s_140_7), .C(CLK_3P3_MHZ_c), .D(n2015));   // src/ram.vhd(56[12:17])
    SB_DFF i3392_3393 (.Q(ram_s_140_6), .C(CLK_3P3_MHZ_c), .D(n2014));   // src/ram.vhd(56[12:17])
    SB_DFF i3389_3390 (.Q(ram_s_140_5), .C(CLK_3P3_MHZ_c), .D(n2013));   // src/ram.vhd(56[12:17])
    SB_DFF i3386_3387 (.Q(ram_s_140_4), .C(CLK_3P3_MHZ_c), .D(n2012));   // src/ram.vhd(56[12:17])
    SB_DFF i3383_3384 (.Q(ram_s_140_3), .C(CLK_3P3_MHZ_c), .D(n2011));   // src/ram.vhd(56[12:17])
    SB_DFF i3380_3381 (.Q(ram_s_140_2), .C(CLK_3P3_MHZ_c), .D(n2010));   // src/ram.vhd(56[12:17])
    SB_DFF i3377_3378 (.Q(ram_s_140_1), .C(CLK_3P3_MHZ_c), .D(n2009));   // src/ram.vhd(56[12:17])
    SB_DFF i3374_3375 (.Q(ram_s_140_0), .C(CLK_3P3_MHZ_c), .D(n2008));   // src/ram.vhd(56[12:17])
    SB_DFF i3371_3372 (.Q(ram_s_139_7), .C(CLK_3P3_MHZ_c), .D(n2007));   // src/ram.vhd(56[12:17])
    SB_DFF i3368_3369 (.Q(ram_s_139_6), .C(CLK_3P3_MHZ_c), .D(n2006));   // src/ram.vhd(56[12:17])
    SB_DFF i3365_3366 (.Q(ram_s_139_5), .C(CLK_3P3_MHZ_c), .D(n2005));   // src/ram.vhd(56[12:17])
    SB_DFF i3362_3363 (.Q(ram_s_139_4), .C(CLK_3P3_MHZ_c), .D(n2004));   // src/ram.vhd(56[12:17])
    SB_DFF i3359_3360 (.Q(ram_s_139_3), .C(CLK_3P3_MHZ_c), .D(n2003));   // src/ram.vhd(56[12:17])
    SB_DFF i3356_3357 (.Q(ram_s_139_2), .C(CLK_3P3_MHZ_c), .D(n2002));   // src/ram.vhd(56[12:17])
    SB_DFF i3353_3354 (.Q(ram_s_139_1), .C(CLK_3P3_MHZ_c), .D(n2001));   // src/ram.vhd(56[12:17])
    SB_DFF i3350_3351 (.Q(ram_s_139_0), .C(CLK_3P3_MHZ_c), .D(n2000));   // src/ram.vhd(56[12:17])
    SB_DFF i3347_3348 (.Q(ram_s_138_7), .C(CLK_3P3_MHZ_c), .D(n1999));   // src/ram.vhd(56[12:17])
    SB_DFF i3344_3345 (.Q(ram_s_138_6), .C(CLK_3P3_MHZ_c), .D(n1998));   // src/ram.vhd(56[12:17])
    SB_DFF i3341_3342 (.Q(ram_s_138_5), .C(CLK_3P3_MHZ_c), .D(n1997));   // src/ram.vhd(56[12:17])
    SB_DFF i3338_3339 (.Q(ram_s_138_4), .C(CLK_3P3_MHZ_c), .D(n1996));   // src/ram.vhd(56[12:17])
    SB_DFF i3335_3336 (.Q(ram_s_138_3), .C(CLK_3P3_MHZ_c), .D(n1995));   // src/ram.vhd(56[12:17])
    SB_DFF i3332_3333 (.Q(ram_s_138_2), .C(CLK_3P3_MHZ_c), .D(n1994));   // src/ram.vhd(56[12:17])
    SB_DFF i3329_3330 (.Q(ram_s_138_1), .C(CLK_3P3_MHZ_c), .D(n1993));   // src/ram.vhd(56[12:17])
    SB_DFF i3326_3327 (.Q(ram_s_138_0), .C(CLK_3P3_MHZ_c), .D(n1992));   // src/ram.vhd(56[12:17])
    SB_DFF i3323_3324 (.Q(ram_s_137_7), .C(CLK_3P3_MHZ_c), .D(n1991));   // src/ram.vhd(56[12:17])
    SB_DFF i3320_3321 (.Q(ram_s_137_6), .C(CLK_3P3_MHZ_c), .D(n1990));   // src/ram.vhd(56[12:17])
    SB_DFF i3317_3318 (.Q(ram_s_137_5), .C(CLK_3P3_MHZ_c), .D(n1989));   // src/ram.vhd(56[12:17])
    SB_DFF i3314_3315 (.Q(ram_s_137_4), .C(CLK_3P3_MHZ_c), .D(n1988));   // src/ram.vhd(56[12:17])
    SB_DFF i3311_3312 (.Q(ram_s_137_3), .C(CLK_3P3_MHZ_c), .D(n1987));   // src/ram.vhd(56[12:17])
    SB_DFF i3308_3309 (.Q(ram_s_137_2), .C(CLK_3P3_MHZ_c), .D(n1986));   // src/ram.vhd(56[12:17])
    SB_DFF i3305_3306 (.Q(ram_s_137_1), .C(CLK_3P3_MHZ_c), .D(n1985));   // src/ram.vhd(56[12:17])
    SB_DFF i3302_3303 (.Q(ram_s_137_0), .C(CLK_3P3_MHZ_c), .D(n1984));   // src/ram.vhd(56[12:17])
    SB_DFF i3299_3300 (.Q(ram_s_136_7), .C(CLK_3P3_MHZ_c), .D(n1983));   // src/ram.vhd(56[12:17])
    SB_DFF i3296_3297 (.Q(ram_s_136_6), .C(CLK_3P3_MHZ_c), .D(n1982));   // src/ram.vhd(56[12:17])
    SB_DFF i3293_3294 (.Q(ram_s_136_5), .C(CLK_3P3_MHZ_c), .D(n1981));   // src/ram.vhd(56[12:17])
    SB_DFF i3290_3291 (.Q(ram_s_136_4), .C(CLK_3P3_MHZ_c), .D(n1980));   // src/ram.vhd(56[12:17])
    SB_DFF i3287_3288 (.Q(ram_s_136_3), .C(CLK_3P3_MHZ_c), .D(n1979));   // src/ram.vhd(56[12:17])
    SB_DFF i3284_3285 (.Q(ram_s_136_2), .C(CLK_3P3_MHZ_c), .D(n1978));   // src/ram.vhd(56[12:17])
    SB_DFF i3281_3282 (.Q(ram_s_136_1), .C(CLK_3P3_MHZ_c), .D(n1977));   // src/ram.vhd(56[12:17])
    SB_DFF i3278_3279 (.Q(ram_s_136_0), .C(CLK_3P3_MHZ_c), .D(n1976));   // src/ram.vhd(56[12:17])
    SB_DFF i3275_3276 (.Q(ram_s_135_7), .C(CLK_3P3_MHZ_c), .D(n1975));   // src/ram.vhd(56[12:17])
    SB_DFF i3272_3273 (.Q(ram_s_135_6), .C(CLK_3P3_MHZ_c), .D(n1974));   // src/ram.vhd(56[12:17])
    SB_DFF i3269_3270 (.Q(ram_s_135_5), .C(CLK_3P3_MHZ_c), .D(n1973));   // src/ram.vhd(56[12:17])
    SB_DFF i3266_3267 (.Q(ram_s_135_4), .C(CLK_3P3_MHZ_c), .D(n1972));   // src/ram.vhd(56[12:17])
    SB_DFF i3263_3264 (.Q(ram_s_135_3), .C(CLK_3P3_MHZ_c), .D(n1971));   // src/ram.vhd(56[12:17])
    SB_DFF i3260_3261 (.Q(ram_s_135_2), .C(CLK_3P3_MHZ_c), .D(n1970));   // src/ram.vhd(56[12:17])
    SB_DFF i3257_3258 (.Q(ram_s_135_1), .C(CLK_3P3_MHZ_c), .D(n1969));   // src/ram.vhd(56[12:17])
    SB_DFF i3254_3255 (.Q(ram_s_135_0), .C(CLK_3P3_MHZ_c), .D(n1968));   // src/ram.vhd(56[12:17])
    SB_DFF i3251_3252 (.Q(ram_s_134_7), .C(CLK_3P3_MHZ_c), .D(n1967));   // src/ram.vhd(56[12:17])
    SB_DFF i3248_3249 (.Q(ram_s_134_6), .C(CLK_3P3_MHZ_c), .D(n1966));   // src/ram.vhd(56[12:17])
    SB_DFF i3245_3246 (.Q(ram_s_134_5), .C(CLK_3P3_MHZ_c), .D(n1965));   // src/ram.vhd(56[12:17])
    SB_DFF i3242_3243 (.Q(ram_s_134_4), .C(CLK_3P3_MHZ_c), .D(n1964));   // src/ram.vhd(56[12:17])
    SB_DFF i3239_3240 (.Q(ram_s_134_3), .C(CLK_3P3_MHZ_c), .D(n1963));   // src/ram.vhd(56[12:17])
    SB_DFF i3236_3237 (.Q(ram_s_134_2), .C(CLK_3P3_MHZ_c), .D(n1962));   // src/ram.vhd(56[12:17])
    SB_DFF i3233_3234 (.Q(ram_s_134_1), .C(CLK_3P3_MHZ_c), .D(n1961));   // src/ram.vhd(56[12:17])
    SB_DFF i3230_3231 (.Q(ram_s_134_0), .C(CLK_3P3_MHZ_c), .D(n1960));   // src/ram.vhd(56[12:17])
    SB_DFF i3227_3228 (.Q(ram_s_133_7), .C(CLK_3P3_MHZ_c), .D(n1959));   // src/ram.vhd(56[12:17])
    SB_DFF i3224_3225 (.Q(ram_s_133_6), .C(CLK_3P3_MHZ_c), .D(n1958));   // src/ram.vhd(56[12:17])
    SB_DFF i3221_3222 (.Q(ram_s_133_5), .C(CLK_3P3_MHZ_c), .D(n1957));   // src/ram.vhd(56[12:17])
    SB_DFF i3218_3219 (.Q(ram_s_133_4), .C(CLK_3P3_MHZ_c), .D(n1956));   // src/ram.vhd(56[12:17])
    SB_DFF i3215_3216 (.Q(ram_s_133_3), .C(CLK_3P3_MHZ_c), .D(n1955));   // src/ram.vhd(56[12:17])
    SB_DFF i3212_3213 (.Q(ram_s_133_2), .C(CLK_3P3_MHZ_c), .D(n1954));   // src/ram.vhd(56[12:17])
    SB_DFF i3209_3210 (.Q(ram_s_133_1), .C(CLK_3P3_MHZ_c), .D(n1953));   // src/ram.vhd(56[12:17])
    SB_DFF i3206_3207 (.Q(ram_s_133_0), .C(CLK_3P3_MHZ_c), .D(n1952));   // src/ram.vhd(56[12:17])
    SB_DFF i3203_3204 (.Q(ram_s_132_7), .C(CLK_3P3_MHZ_c), .D(n1951));   // src/ram.vhd(56[12:17])
    SB_DFF i3200_3201 (.Q(ram_s_132_6), .C(CLK_3P3_MHZ_c), .D(n1950));   // src/ram.vhd(56[12:17])
    SB_DFF i3197_3198 (.Q(ram_s_132_5), .C(CLK_3P3_MHZ_c), .D(n1949));   // src/ram.vhd(56[12:17])
    SB_DFF i3194_3195 (.Q(ram_s_132_4), .C(CLK_3P3_MHZ_c), .D(n1948));   // src/ram.vhd(56[12:17])
    SB_DFF i3191_3192 (.Q(ram_s_132_3), .C(CLK_3P3_MHZ_c), .D(n1947));   // src/ram.vhd(56[12:17])
    SB_DFF i3188_3189 (.Q(ram_s_132_2), .C(CLK_3P3_MHZ_c), .D(n1946));   // src/ram.vhd(56[12:17])
    SB_DFF i3185_3186 (.Q(ram_s_132_1), .C(CLK_3P3_MHZ_c), .D(n1945));   // src/ram.vhd(56[12:17])
    SB_DFF i3182_3183 (.Q(ram_s_132_0), .C(CLK_3P3_MHZ_c), .D(n1944));   // src/ram.vhd(56[12:17])
    SB_DFF i3179_3180 (.Q(ram_s_131_7), .C(CLK_3P3_MHZ_c), .D(n1943));   // src/ram.vhd(56[12:17])
    SB_DFF i3176_3177 (.Q(ram_s_131_6), .C(CLK_3P3_MHZ_c), .D(n1942));   // src/ram.vhd(56[12:17])
    SB_DFF i3173_3174 (.Q(ram_s_131_5), .C(CLK_3P3_MHZ_c), .D(n1941));   // src/ram.vhd(56[12:17])
    SB_DFF i3170_3171 (.Q(ram_s_131_4), .C(CLK_3P3_MHZ_c), .D(n1940));   // src/ram.vhd(56[12:17])
    SB_DFF i3167_3168 (.Q(ram_s_131_3), .C(CLK_3P3_MHZ_c), .D(n1939));   // src/ram.vhd(56[12:17])
    SB_DFF i3164_3165 (.Q(ram_s_131_2), .C(CLK_3P3_MHZ_c), .D(n1938));   // src/ram.vhd(56[12:17])
    SB_DFF i3161_3162 (.Q(ram_s_131_1), .C(CLK_3P3_MHZ_c), .D(n1937));   // src/ram.vhd(56[12:17])
    SB_DFF i3158_3159 (.Q(ram_s_131_0), .C(CLK_3P3_MHZ_c), .D(n1936));   // src/ram.vhd(56[12:17])
    SB_DFF i3155_3156 (.Q(ram_s_130_7), .C(CLK_3P3_MHZ_c), .D(n1935));   // src/ram.vhd(56[12:17])
    SB_DFF i3152_3153 (.Q(ram_s_130_6), .C(CLK_3P3_MHZ_c), .D(n1934));   // src/ram.vhd(56[12:17])
    SB_DFF i3149_3150 (.Q(ram_s_130_5), .C(CLK_3P3_MHZ_c), .D(n1933));   // src/ram.vhd(56[12:17])
    SB_DFF i3146_3147 (.Q(ram_s_130_4), .C(CLK_3P3_MHZ_c), .D(n1932));   // src/ram.vhd(56[12:17])
    SB_DFF i3143_3144 (.Q(ram_s_130_3), .C(CLK_3P3_MHZ_c), .D(n1931));   // src/ram.vhd(56[12:17])
    SB_DFF i3140_3141 (.Q(ram_s_130_2), .C(CLK_3P3_MHZ_c), .D(n1930));   // src/ram.vhd(56[12:17])
    SB_DFF i3137_3138 (.Q(ram_s_130_1), .C(CLK_3P3_MHZ_c), .D(n1929));   // src/ram.vhd(56[12:17])
    SB_DFF i3134_3135 (.Q(ram_s_130_0), .C(CLK_3P3_MHZ_c), .D(n1928));   // src/ram.vhd(56[12:17])
    SB_DFF i3131_3132 (.Q(ram_s_129_7), .C(CLK_3P3_MHZ_c), .D(n1927));   // src/ram.vhd(56[12:17])
    SB_DFF i3128_3129 (.Q(ram_s_129_6), .C(CLK_3P3_MHZ_c), .D(n1926));   // src/ram.vhd(56[12:17])
    SB_DFF i3125_3126 (.Q(ram_s_129_5), .C(CLK_3P3_MHZ_c), .D(n1925));   // src/ram.vhd(56[12:17])
    SB_DFF i3122_3123 (.Q(ram_s_129_4), .C(CLK_3P3_MHZ_c), .D(n1924));   // src/ram.vhd(56[12:17])
    SB_DFF i3119_3120 (.Q(ram_s_129_3), .C(CLK_3P3_MHZ_c), .D(n1923));   // src/ram.vhd(56[12:17])
    SB_DFF i3116_3117 (.Q(ram_s_129_2), .C(CLK_3P3_MHZ_c), .D(n1922));   // src/ram.vhd(56[12:17])
    SB_DFF i3113_3114 (.Q(ram_s_129_1), .C(CLK_3P3_MHZ_c), .D(n1921));   // src/ram.vhd(56[12:17])
    SB_DFF i3110_3111 (.Q(ram_s_129_0), .C(CLK_3P3_MHZ_c), .D(n1920));   // src/ram.vhd(56[12:17])
    SB_DFF i3107_3108 (.Q(ram_s_128_7), .C(CLK_3P3_MHZ_c), .D(n1919));   // src/ram.vhd(56[12:17])
    SB_DFF i3104_3105 (.Q(ram_s_128_6), .C(CLK_3P3_MHZ_c), .D(n1918));   // src/ram.vhd(56[12:17])
    SB_DFF i3101_3102 (.Q(ram_s_128_5), .C(CLK_3P3_MHZ_c), .D(n1917));   // src/ram.vhd(56[12:17])
    SB_DFF i3098_3099 (.Q(ram_s_128_4), .C(CLK_3P3_MHZ_c), .D(n1916));   // src/ram.vhd(56[12:17])
    SB_DFF i3095_3096 (.Q(ram_s_128_3), .C(CLK_3P3_MHZ_c), .D(n1915));   // src/ram.vhd(56[12:17])
    SB_DFF i3092_3093 (.Q(ram_s_128_2), .C(CLK_3P3_MHZ_c), .D(n1914));   // src/ram.vhd(56[12:17])
    SB_DFF i3089_3090 (.Q(ram_s_128_1), .C(CLK_3P3_MHZ_c), .D(n1913));   // src/ram.vhd(56[12:17])
    SB_DFF i3086_3087 (.Q(ram_s_128_0), .C(CLK_3P3_MHZ_c), .D(n1912));   // src/ram.vhd(56[12:17])
    SB_DFF i3083_3084 (.Q(ram_s_127_7), .C(CLK_3P3_MHZ_c), .D(n1911));   // src/ram.vhd(56[12:17])
    SB_DFF i3080_3081 (.Q(ram_s_127_6), .C(CLK_3P3_MHZ_c), .D(n1910));   // src/ram.vhd(56[12:17])
    SB_DFF i3077_3078 (.Q(ram_s_127_5), .C(CLK_3P3_MHZ_c), .D(n1909));   // src/ram.vhd(56[12:17])
    SB_DFF i3074_3075 (.Q(ram_s_127_4), .C(CLK_3P3_MHZ_c), .D(n1908));   // src/ram.vhd(56[12:17])
    SB_DFF i3071_3072 (.Q(ram_s_127_3), .C(CLK_3P3_MHZ_c), .D(n1907));   // src/ram.vhd(56[12:17])
    SB_DFF i3068_3069 (.Q(ram_s_127_2), .C(CLK_3P3_MHZ_c), .D(n1906));   // src/ram.vhd(56[12:17])
    SB_DFF i3065_3066 (.Q(ram_s_127_1), .C(CLK_3P3_MHZ_c), .D(n1905));   // src/ram.vhd(56[12:17])
    SB_DFF i3062_3063 (.Q(ram_s_127_0), .C(CLK_3P3_MHZ_c), .D(n1904));   // src/ram.vhd(56[12:17])
    SB_DFF i3059_3060 (.Q(ram_s_126_7), .C(CLK_3P3_MHZ_c), .D(n1903));   // src/ram.vhd(56[12:17])
    SB_DFF i3056_3057 (.Q(ram_s_126_6), .C(CLK_3P3_MHZ_c), .D(n1902));   // src/ram.vhd(56[12:17])
    SB_DFF i3053_3054 (.Q(ram_s_126_5), .C(CLK_3P3_MHZ_c), .D(n1901));   // src/ram.vhd(56[12:17])
    SB_DFF i3050_3051 (.Q(ram_s_126_4), .C(CLK_3P3_MHZ_c), .D(n1900));   // src/ram.vhd(56[12:17])
    SB_DFF i3047_3048 (.Q(ram_s_126_3), .C(CLK_3P3_MHZ_c), .D(n1899));   // src/ram.vhd(56[12:17])
    SB_DFF i3044_3045 (.Q(ram_s_126_2), .C(CLK_3P3_MHZ_c), .D(n1898));   // src/ram.vhd(56[12:17])
    SB_DFF i3041_3042 (.Q(ram_s_126_1), .C(CLK_3P3_MHZ_c), .D(n1897));   // src/ram.vhd(56[12:17])
    SB_DFF i3038_3039 (.Q(ram_s_126_0), .C(CLK_3P3_MHZ_c), .D(n1896));   // src/ram.vhd(56[12:17])
    SB_DFF i3035_3036 (.Q(ram_s_125_7), .C(CLK_3P3_MHZ_c), .D(n1895));   // src/ram.vhd(56[12:17])
    SB_DFF i3032_3033 (.Q(ram_s_125_6), .C(CLK_3P3_MHZ_c), .D(n1894));   // src/ram.vhd(56[12:17])
    SB_DFF i3029_3030 (.Q(ram_s_125_5), .C(CLK_3P3_MHZ_c), .D(n1893));   // src/ram.vhd(56[12:17])
    SB_DFF i3026_3027 (.Q(ram_s_125_4), .C(CLK_3P3_MHZ_c), .D(n1892));   // src/ram.vhd(56[12:17])
    SB_DFF i3023_3024 (.Q(ram_s_125_3), .C(CLK_3P3_MHZ_c), .D(n1891));   // src/ram.vhd(56[12:17])
    SB_DFF i3020_3021 (.Q(ram_s_125_2), .C(CLK_3P3_MHZ_c), .D(n1890));   // src/ram.vhd(56[12:17])
    SB_DFF i3017_3018 (.Q(ram_s_125_1), .C(CLK_3P3_MHZ_c), .D(n1889));   // src/ram.vhd(56[12:17])
    SB_DFF i3014_3015 (.Q(ram_s_125_0), .C(CLK_3P3_MHZ_c), .D(n1888));   // src/ram.vhd(56[12:17])
    SB_DFF i3011_3012 (.Q(ram_s_124_7), .C(CLK_3P3_MHZ_c), .D(n1887));   // src/ram.vhd(56[12:17])
    SB_DFF i3008_3009 (.Q(ram_s_124_6), .C(CLK_3P3_MHZ_c), .D(n1886));   // src/ram.vhd(56[12:17])
    SB_DFF i3005_3006 (.Q(ram_s_124_5), .C(CLK_3P3_MHZ_c), .D(n1885));   // src/ram.vhd(56[12:17])
    SB_DFF i3002_3003 (.Q(ram_s_124_4), .C(CLK_3P3_MHZ_c), .D(n1884));   // src/ram.vhd(56[12:17])
    SB_DFF i2999_3000 (.Q(ram_s_124_3), .C(CLK_3P3_MHZ_c), .D(n1883));   // src/ram.vhd(56[12:17])
    SB_DFF i2996_2997 (.Q(ram_s_124_2), .C(CLK_3P3_MHZ_c), .D(n1882));   // src/ram.vhd(56[12:17])
    SB_DFF i2993_2994 (.Q(ram_s_124_1), .C(CLK_3P3_MHZ_c), .D(n1881));   // src/ram.vhd(56[12:17])
    SB_DFF i2990_2991 (.Q(ram_s_124_0), .C(CLK_3P3_MHZ_c), .D(n1880));   // src/ram.vhd(56[12:17])
    SB_DFF i2987_2988 (.Q(ram_s_123_7), .C(CLK_3P3_MHZ_c), .D(n1879));   // src/ram.vhd(56[12:17])
    SB_DFF i2984_2985 (.Q(ram_s_123_6), .C(CLK_3P3_MHZ_c), .D(n1878));   // src/ram.vhd(56[12:17])
    SB_DFF i2981_2982 (.Q(ram_s_123_5), .C(CLK_3P3_MHZ_c), .D(n1877));   // src/ram.vhd(56[12:17])
    SB_DFF i2978_2979 (.Q(ram_s_123_4), .C(CLK_3P3_MHZ_c), .D(n1876));   // src/ram.vhd(56[12:17])
    SB_DFF i2975_2976 (.Q(ram_s_123_3), .C(CLK_3P3_MHZ_c), .D(n1875));   // src/ram.vhd(56[12:17])
    SB_DFF i2972_2973 (.Q(ram_s_123_2), .C(CLK_3P3_MHZ_c), .D(n1874));   // src/ram.vhd(56[12:17])
    SB_DFF i2969_2970 (.Q(ram_s_123_1), .C(CLK_3P3_MHZ_c), .D(n1873));   // src/ram.vhd(56[12:17])
    SB_DFF i2966_2967 (.Q(ram_s_123_0), .C(CLK_3P3_MHZ_c), .D(n1872));   // src/ram.vhd(56[12:17])
    SB_DFF i2963_2964 (.Q(ram_s_122_7), .C(CLK_3P3_MHZ_c), .D(n1871));   // src/ram.vhd(56[12:17])
    SB_DFF i2960_2961 (.Q(ram_s_122_6), .C(CLK_3P3_MHZ_c), .D(n1870));   // src/ram.vhd(56[12:17])
    SB_DFF i2957_2958 (.Q(ram_s_122_5), .C(CLK_3P3_MHZ_c), .D(n1869));   // src/ram.vhd(56[12:17])
    SB_DFF i2954_2955 (.Q(ram_s_122_4), .C(CLK_3P3_MHZ_c), .D(n1868));   // src/ram.vhd(56[12:17])
    SB_DFF i2951_2952 (.Q(ram_s_122_3), .C(CLK_3P3_MHZ_c), .D(n1867));   // src/ram.vhd(56[12:17])
    SB_DFF i2948_2949 (.Q(ram_s_122_2), .C(CLK_3P3_MHZ_c), .D(n1866));   // src/ram.vhd(56[12:17])
    SB_DFF i2945_2946 (.Q(ram_s_122_1), .C(CLK_3P3_MHZ_c), .D(n1865));   // src/ram.vhd(56[12:17])
    SB_DFF i2942_2943 (.Q(ram_s_122_0), .C(CLK_3P3_MHZ_c), .D(n1864));   // src/ram.vhd(56[12:17])
    SB_DFF i2939_2940 (.Q(ram_s_121_7), .C(CLK_3P3_MHZ_c), .D(n1863));   // src/ram.vhd(56[12:17])
    SB_DFF i2936_2937 (.Q(ram_s_121_6), .C(CLK_3P3_MHZ_c), .D(n1862));   // src/ram.vhd(56[12:17])
    SB_DFF i2933_2934 (.Q(ram_s_121_5), .C(CLK_3P3_MHZ_c), .D(n1861));   // src/ram.vhd(56[12:17])
    SB_DFF i2930_2931 (.Q(ram_s_121_4), .C(CLK_3P3_MHZ_c), .D(n1860));   // src/ram.vhd(56[12:17])
    SB_DFF i2927_2928 (.Q(ram_s_121_3), .C(CLK_3P3_MHZ_c), .D(n1859));   // src/ram.vhd(56[12:17])
    SB_DFF i2924_2925 (.Q(ram_s_121_2), .C(CLK_3P3_MHZ_c), .D(n1858));   // src/ram.vhd(56[12:17])
    SB_DFF i2921_2922 (.Q(ram_s_121_1), .C(CLK_3P3_MHZ_c), .D(n1857));   // src/ram.vhd(56[12:17])
    SB_DFF i2918_2919 (.Q(ram_s_121_0), .C(CLK_3P3_MHZ_c), .D(n1856));   // src/ram.vhd(56[12:17])
    SB_DFF i2915_2916 (.Q(ram_s_120_7), .C(CLK_3P3_MHZ_c), .D(n1855));   // src/ram.vhd(56[12:17])
    SB_DFF i2912_2913 (.Q(ram_s_120_6), .C(CLK_3P3_MHZ_c), .D(n1854));   // src/ram.vhd(56[12:17])
    SB_DFF i2909_2910 (.Q(ram_s_120_5), .C(CLK_3P3_MHZ_c), .D(n1853));   // src/ram.vhd(56[12:17])
    SB_DFF i2906_2907 (.Q(ram_s_120_4), .C(CLK_3P3_MHZ_c), .D(n1852));   // src/ram.vhd(56[12:17])
    SB_DFF i2903_2904 (.Q(ram_s_120_3), .C(CLK_3P3_MHZ_c), .D(n1851));   // src/ram.vhd(56[12:17])
    SB_DFF i2900_2901 (.Q(ram_s_120_2), .C(CLK_3P3_MHZ_c), .D(n1850));   // src/ram.vhd(56[12:17])
    SB_DFF i2897_2898 (.Q(ram_s_120_1), .C(CLK_3P3_MHZ_c), .D(n1849));   // src/ram.vhd(56[12:17])
    SB_DFF i2894_2895 (.Q(ram_s_120_0), .C(CLK_3P3_MHZ_c), .D(n1848));   // src/ram.vhd(56[12:17])
    SB_DFF i2891_2892 (.Q(ram_s_119_7), .C(CLK_3P3_MHZ_c), .D(n1847));   // src/ram.vhd(56[12:17])
    SB_DFF i2888_2889 (.Q(ram_s_119_6), .C(CLK_3P3_MHZ_c), .D(n1846));   // src/ram.vhd(56[12:17])
    SB_DFF i2885_2886 (.Q(ram_s_119_5), .C(CLK_3P3_MHZ_c), .D(n1845));   // src/ram.vhd(56[12:17])
    SB_DFF i2882_2883 (.Q(ram_s_119_4), .C(CLK_3P3_MHZ_c), .D(n1844));   // src/ram.vhd(56[12:17])
    SB_DFF i2879_2880 (.Q(ram_s_119_3), .C(CLK_3P3_MHZ_c), .D(n1843));   // src/ram.vhd(56[12:17])
    SB_DFF i2876_2877 (.Q(ram_s_119_2), .C(CLK_3P3_MHZ_c), .D(n1842));   // src/ram.vhd(56[12:17])
    SB_DFF i2873_2874 (.Q(ram_s_119_1), .C(CLK_3P3_MHZ_c), .D(n1841));   // src/ram.vhd(56[12:17])
    SB_DFF i2870_2871 (.Q(ram_s_119_0), .C(CLK_3P3_MHZ_c), .D(n1840));   // src/ram.vhd(56[12:17])
    SB_DFF i2867_2868 (.Q(ram_s_118_7), .C(CLK_3P3_MHZ_c), .D(n1839));   // src/ram.vhd(56[12:17])
    SB_DFF i2864_2865 (.Q(ram_s_118_6), .C(CLK_3P3_MHZ_c), .D(n1838));   // src/ram.vhd(56[12:17])
    SB_DFF i2861_2862 (.Q(ram_s_118_5), .C(CLK_3P3_MHZ_c), .D(n1837));   // src/ram.vhd(56[12:17])
    SB_DFF i2858_2859 (.Q(ram_s_118_4), .C(CLK_3P3_MHZ_c), .D(n1836));   // src/ram.vhd(56[12:17])
    SB_DFF i2855_2856 (.Q(ram_s_118_3), .C(CLK_3P3_MHZ_c), .D(n1835));   // src/ram.vhd(56[12:17])
    SB_DFF i2852_2853 (.Q(ram_s_118_2), .C(CLK_3P3_MHZ_c), .D(n1834));   // src/ram.vhd(56[12:17])
    SB_DFF i2849_2850 (.Q(ram_s_118_1), .C(CLK_3P3_MHZ_c), .D(n1833));   // src/ram.vhd(56[12:17])
    SB_DFF i2846_2847 (.Q(ram_s_118_0), .C(CLK_3P3_MHZ_c), .D(n1832));   // src/ram.vhd(56[12:17])
    SB_DFF i2843_2844 (.Q(ram_s_117_7), .C(CLK_3P3_MHZ_c), .D(n1831));   // src/ram.vhd(56[12:17])
    SB_DFF i2840_2841 (.Q(ram_s_117_6), .C(CLK_3P3_MHZ_c), .D(n1830));   // src/ram.vhd(56[12:17])
    SB_DFF i2837_2838 (.Q(ram_s_117_5), .C(CLK_3P3_MHZ_c), .D(n1829));   // src/ram.vhd(56[12:17])
    SB_DFF i2834_2835 (.Q(ram_s_117_4), .C(CLK_3P3_MHZ_c), .D(n1828));   // src/ram.vhd(56[12:17])
    SB_DFF i2831_2832 (.Q(ram_s_117_3), .C(CLK_3P3_MHZ_c), .D(n1827));   // src/ram.vhd(56[12:17])
    SB_DFF i2828_2829 (.Q(ram_s_117_2), .C(CLK_3P3_MHZ_c), .D(n1826));   // src/ram.vhd(56[12:17])
    SB_DFF i2825_2826 (.Q(ram_s_117_1), .C(CLK_3P3_MHZ_c), .D(n1825));   // src/ram.vhd(56[12:17])
    SB_DFF i2822_2823 (.Q(ram_s_117_0), .C(CLK_3P3_MHZ_c), .D(n1824));   // src/ram.vhd(56[12:17])
    SB_DFF i2819_2820 (.Q(ram_s_116_7), .C(CLK_3P3_MHZ_c), .D(n1823));   // src/ram.vhd(56[12:17])
    SB_DFF i2816_2817 (.Q(ram_s_116_6), .C(CLK_3P3_MHZ_c), .D(n1822));   // src/ram.vhd(56[12:17])
    SB_DFF i2813_2814 (.Q(ram_s_116_5), .C(CLK_3P3_MHZ_c), .D(n1821));   // src/ram.vhd(56[12:17])
    SB_DFF i2810_2811 (.Q(ram_s_116_4), .C(CLK_3P3_MHZ_c), .D(n1820));   // src/ram.vhd(56[12:17])
    SB_DFF i2807_2808 (.Q(ram_s_116_3), .C(CLK_3P3_MHZ_c), .D(n1819));   // src/ram.vhd(56[12:17])
    SB_DFF i2804_2805 (.Q(ram_s_116_2), .C(CLK_3P3_MHZ_c), .D(n1818));   // src/ram.vhd(56[12:17])
    SB_DFF i2801_2802 (.Q(ram_s_116_1), .C(CLK_3P3_MHZ_c), .D(n1817));   // src/ram.vhd(56[12:17])
    SB_DFF i2798_2799 (.Q(ram_s_116_0), .C(CLK_3P3_MHZ_c), .D(n1816));   // src/ram.vhd(56[12:17])
    SB_DFF i2795_2796 (.Q(ram_s_115_7), .C(CLK_3P3_MHZ_c), .D(n1815));   // src/ram.vhd(56[12:17])
    SB_DFF i2792_2793 (.Q(ram_s_115_6), .C(CLK_3P3_MHZ_c), .D(n1814));   // src/ram.vhd(56[12:17])
    SB_DFF i2789_2790 (.Q(ram_s_115_5), .C(CLK_3P3_MHZ_c), .D(n1813));   // src/ram.vhd(56[12:17])
    SB_DFF i2786_2787 (.Q(ram_s_115_4), .C(CLK_3P3_MHZ_c), .D(n1812));   // src/ram.vhd(56[12:17])
    SB_DFF i2783_2784 (.Q(ram_s_115_3), .C(CLK_3P3_MHZ_c), .D(n1811));   // src/ram.vhd(56[12:17])
    SB_DFF i2780_2781 (.Q(ram_s_115_2), .C(CLK_3P3_MHZ_c), .D(n1810));   // src/ram.vhd(56[12:17])
    SB_DFF i2777_2778 (.Q(ram_s_115_1), .C(CLK_3P3_MHZ_c), .D(n1809));   // src/ram.vhd(56[12:17])
    SB_DFF i2774_2775 (.Q(ram_s_115_0), .C(CLK_3P3_MHZ_c), .D(n1808));   // src/ram.vhd(56[12:17])
    SB_DFF i2771_2772 (.Q(ram_s_114_7), .C(CLK_3P3_MHZ_c), .D(n1807));   // src/ram.vhd(56[12:17])
    SB_DFF i2768_2769 (.Q(ram_s_114_6), .C(CLK_3P3_MHZ_c), .D(n1806));   // src/ram.vhd(56[12:17])
    SB_DFF i2765_2766 (.Q(ram_s_114_5), .C(CLK_3P3_MHZ_c), .D(n1805));   // src/ram.vhd(56[12:17])
    SB_DFF i2762_2763 (.Q(ram_s_114_4), .C(CLK_3P3_MHZ_c), .D(n1804));   // src/ram.vhd(56[12:17])
    SB_DFF i2759_2760 (.Q(ram_s_114_3), .C(CLK_3P3_MHZ_c), .D(n1803));   // src/ram.vhd(56[12:17])
    SB_DFF i2756_2757 (.Q(ram_s_114_2), .C(CLK_3P3_MHZ_c), .D(n1802));   // src/ram.vhd(56[12:17])
    SB_DFF i2753_2754 (.Q(ram_s_114_1), .C(CLK_3P3_MHZ_c), .D(n1801));   // src/ram.vhd(56[12:17])
    SB_DFF i2750_2751 (.Q(ram_s_114_0), .C(CLK_3P3_MHZ_c), .D(n1800));   // src/ram.vhd(56[12:17])
    SB_DFF i2747_2748 (.Q(ram_s_113_7), .C(CLK_3P3_MHZ_c), .D(n1799));   // src/ram.vhd(56[12:17])
    SB_DFF i2744_2745 (.Q(ram_s_113_6), .C(CLK_3P3_MHZ_c), .D(n1798));   // src/ram.vhd(56[12:17])
    SB_DFF i2741_2742 (.Q(ram_s_113_5), .C(CLK_3P3_MHZ_c), .D(n1797));   // src/ram.vhd(56[12:17])
    SB_DFF i2738_2739 (.Q(ram_s_113_4), .C(CLK_3P3_MHZ_c), .D(n1796));   // src/ram.vhd(56[12:17])
    SB_DFF i2735_2736 (.Q(ram_s_113_3), .C(CLK_3P3_MHZ_c), .D(n1795));   // src/ram.vhd(56[12:17])
    SB_DFF i2732_2733 (.Q(ram_s_113_2), .C(CLK_3P3_MHZ_c), .D(n1794));   // src/ram.vhd(56[12:17])
    SB_DFF i2729_2730 (.Q(ram_s_113_1), .C(CLK_3P3_MHZ_c), .D(n1793));   // src/ram.vhd(56[12:17])
    SB_DFF i2726_2727 (.Q(ram_s_113_0), .C(CLK_3P3_MHZ_c), .D(n1792));   // src/ram.vhd(56[12:17])
    SB_DFF i2723_2724 (.Q(ram_s_112_7), .C(CLK_3P3_MHZ_c), .D(n1791));   // src/ram.vhd(56[12:17])
    SB_DFF i2720_2721 (.Q(ram_s_112_6), .C(CLK_3P3_MHZ_c), .D(n1790));   // src/ram.vhd(56[12:17])
    SB_DFF i2717_2718 (.Q(ram_s_112_5), .C(CLK_3P3_MHZ_c), .D(n1789));   // src/ram.vhd(56[12:17])
    SB_DFF i2714_2715 (.Q(ram_s_112_4), .C(CLK_3P3_MHZ_c), .D(n1788));   // src/ram.vhd(56[12:17])
    SB_DFF i2711_2712 (.Q(ram_s_112_3), .C(CLK_3P3_MHZ_c), .D(n1787));   // src/ram.vhd(56[12:17])
    SB_DFF i2708_2709 (.Q(ram_s_112_2), .C(CLK_3P3_MHZ_c), .D(n1786));   // src/ram.vhd(56[12:17])
    SB_DFF i2705_2706 (.Q(ram_s_112_1), .C(CLK_3P3_MHZ_c), .D(n1785));   // src/ram.vhd(56[12:17])
    SB_DFF i2702_2703 (.Q(ram_s_112_0), .C(CLK_3P3_MHZ_c), .D(n1784));   // src/ram.vhd(56[12:17])
    SB_DFF i2699_2700 (.Q(ram_s_111_7), .C(CLK_3P3_MHZ_c), .D(n1783));   // src/ram.vhd(56[12:17])
    SB_DFF i2696_2697 (.Q(ram_s_111_6), .C(CLK_3P3_MHZ_c), .D(n1782));   // src/ram.vhd(56[12:17])
    SB_DFF i2693_2694 (.Q(ram_s_111_5), .C(CLK_3P3_MHZ_c), .D(n1781));   // src/ram.vhd(56[12:17])
    SB_DFF i2690_2691 (.Q(ram_s_111_4), .C(CLK_3P3_MHZ_c), .D(n1780));   // src/ram.vhd(56[12:17])
    SB_DFF i2687_2688 (.Q(ram_s_111_3), .C(CLK_3P3_MHZ_c), .D(n1779));   // src/ram.vhd(56[12:17])
    SB_DFF i2684_2685 (.Q(ram_s_111_2), .C(CLK_3P3_MHZ_c), .D(n1778));   // src/ram.vhd(56[12:17])
    SB_DFF i2681_2682 (.Q(ram_s_111_1), .C(CLK_3P3_MHZ_c), .D(n1777));   // src/ram.vhd(56[12:17])
    SB_DFF i2678_2679 (.Q(ram_s_111_0), .C(CLK_3P3_MHZ_c), .D(n1776));   // src/ram.vhd(56[12:17])
    SB_DFF i2675_2676 (.Q(ram_s_110_7), .C(CLK_3P3_MHZ_c), .D(n1775));   // src/ram.vhd(56[12:17])
    SB_DFF i2672_2673 (.Q(ram_s_110_6), .C(CLK_3P3_MHZ_c), .D(n1774));   // src/ram.vhd(56[12:17])
    SB_DFF i2669_2670 (.Q(ram_s_110_5), .C(CLK_3P3_MHZ_c), .D(n1773));   // src/ram.vhd(56[12:17])
    SB_DFF i2666_2667 (.Q(ram_s_110_4), .C(CLK_3P3_MHZ_c), .D(n1772));   // src/ram.vhd(56[12:17])
    SB_DFF i2663_2664 (.Q(ram_s_110_3), .C(CLK_3P3_MHZ_c), .D(n1771));   // src/ram.vhd(56[12:17])
    SB_DFF i2660_2661 (.Q(ram_s_110_2), .C(CLK_3P3_MHZ_c), .D(n1770));   // src/ram.vhd(56[12:17])
    SB_DFF i2657_2658 (.Q(ram_s_110_1), .C(CLK_3P3_MHZ_c), .D(n1769));   // src/ram.vhd(56[12:17])
    SB_DFF i2654_2655 (.Q(ram_s_110_0), .C(CLK_3P3_MHZ_c), .D(n1768));   // src/ram.vhd(56[12:17])
    SB_DFF i2651_2652 (.Q(ram_s_109_7), .C(CLK_3P3_MHZ_c), .D(n1767));   // src/ram.vhd(56[12:17])
    SB_DFF i2648_2649 (.Q(ram_s_109_6), .C(CLK_3P3_MHZ_c), .D(n1766));   // src/ram.vhd(56[12:17])
    SB_DFF i2645_2646 (.Q(ram_s_109_5), .C(CLK_3P3_MHZ_c), .D(n1765));   // src/ram.vhd(56[12:17])
    SB_DFF i2642_2643 (.Q(ram_s_109_4), .C(CLK_3P3_MHZ_c), .D(n1764));   // src/ram.vhd(56[12:17])
    SB_DFF i2639_2640 (.Q(ram_s_109_3), .C(CLK_3P3_MHZ_c), .D(n1763));   // src/ram.vhd(56[12:17])
    SB_DFF i2636_2637 (.Q(ram_s_109_2), .C(CLK_3P3_MHZ_c), .D(n1762));   // src/ram.vhd(56[12:17])
    SB_DFF i2633_2634 (.Q(ram_s_109_1), .C(CLK_3P3_MHZ_c), .D(n1761));   // src/ram.vhd(56[12:17])
    SB_DFF i2630_2631 (.Q(ram_s_109_0), .C(CLK_3P3_MHZ_c), .D(n1760));   // src/ram.vhd(56[12:17])
    SB_DFF i2627_2628 (.Q(ram_s_108_7), .C(CLK_3P3_MHZ_c), .D(n1759));   // src/ram.vhd(56[12:17])
    SB_DFF i2624_2625 (.Q(ram_s_108_6), .C(CLK_3P3_MHZ_c), .D(n1758));   // src/ram.vhd(56[12:17])
    SB_DFF i2621_2622 (.Q(ram_s_108_5), .C(CLK_3P3_MHZ_c), .D(n1757));   // src/ram.vhd(56[12:17])
    SB_DFF i2618_2619 (.Q(ram_s_108_4), .C(CLK_3P3_MHZ_c), .D(n1756));   // src/ram.vhd(56[12:17])
    SB_DFF i2615_2616 (.Q(ram_s_108_3), .C(CLK_3P3_MHZ_c), .D(n1755));   // src/ram.vhd(56[12:17])
    SB_DFF i2612_2613 (.Q(ram_s_108_2), .C(CLK_3P3_MHZ_c), .D(n1754));   // src/ram.vhd(56[12:17])
    SB_DFF i2609_2610 (.Q(ram_s_108_1), .C(CLK_3P3_MHZ_c), .D(n1753));   // src/ram.vhd(56[12:17])
    SB_DFF i2606_2607 (.Q(ram_s_108_0), .C(CLK_3P3_MHZ_c), .D(n1752));   // src/ram.vhd(56[12:17])
    SB_DFF i2603_2604 (.Q(ram_s_107_7), .C(CLK_3P3_MHZ_c), .D(n1751));   // src/ram.vhd(56[12:17])
    SB_DFF i2600_2601 (.Q(ram_s_107_6), .C(CLK_3P3_MHZ_c), .D(n1750));   // src/ram.vhd(56[12:17])
    SB_DFF i2597_2598 (.Q(ram_s_107_5), .C(CLK_3P3_MHZ_c), .D(n1749));   // src/ram.vhd(56[12:17])
    SB_DFF i2594_2595 (.Q(ram_s_107_4), .C(CLK_3P3_MHZ_c), .D(n1748));   // src/ram.vhd(56[12:17])
    SB_DFF i2591_2592 (.Q(ram_s_107_3), .C(CLK_3P3_MHZ_c), .D(n1747));   // src/ram.vhd(56[12:17])
    SB_DFF i2588_2589 (.Q(ram_s_107_2), .C(CLK_3P3_MHZ_c), .D(n1746));   // src/ram.vhd(56[12:17])
    SB_DFF i2585_2586 (.Q(ram_s_107_1), .C(CLK_3P3_MHZ_c), .D(n1745));   // src/ram.vhd(56[12:17])
    SB_DFF i2582_2583 (.Q(ram_s_107_0), .C(CLK_3P3_MHZ_c), .D(n1744));   // src/ram.vhd(56[12:17])
    SB_DFF i2579_2580 (.Q(ram_s_106_7), .C(CLK_3P3_MHZ_c), .D(n1743));   // src/ram.vhd(56[12:17])
    SB_DFF i2576_2577 (.Q(ram_s_106_6), .C(CLK_3P3_MHZ_c), .D(n1742));   // src/ram.vhd(56[12:17])
    SB_DFF i2573_2574 (.Q(ram_s_106_5), .C(CLK_3P3_MHZ_c), .D(n1741));   // src/ram.vhd(56[12:17])
    SB_DFF i2570_2571 (.Q(ram_s_106_4), .C(CLK_3P3_MHZ_c), .D(n1740));   // src/ram.vhd(56[12:17])
    SB_DFF i2567_2568 (.Q(ram_s_106_3), .C(CLK_3P3_MHZ_c), .D(n1739));   // src/ram.vhd(56[12:17])
    SB_DFF i2564_2565 (.Q(ram_s_106_2), .C(CLK_3P3_MHZ_c), .D(n1738));   // src/ram.vhd(56[12:17])
    SB_DFF i2561_2562 (.Q(ram_s_106_1), .C(CLK_3P3_MHZ_c), .D(n1737));   // src/ram.vhd(56[12:17])
    SB_DFF i2558_2559 (.Q(ram_s_106_0), .C(CLK_3P3_MHZ_c), .D(n1736));   // src/ram.vhd(56[12:17])
    SB_DFF i2555_2556 (.Q(ram_s_105_7), .C(CLK_3P3_MHZ_c), .D(n1735));   // src/ram.vhd(56[12:17])
    SB_DFF i2552_2553 (.Q(ram_s_105_6), .C(CLK_3P3_MHZ_c), .D(n1734));   // src/ram.vhd(56[12:17])
    SB_DFF i2549_2550 (.Q(ram_s_105_5), .C(CLK_3P3_MHZ_c), .D(n1733));   // src/ram.vhd(56[12:17])
    SB_DFF i2546_2547 (.Q(ram_s_105_4), .C(CLK_3P3_MHZ_c), .D(n1732));   // src/ram.vhd(56[12:17])
    SB_DFF i2543_2544 (.Q(ram_s_105_3), .C(CLK_3P3_MHZ_c), .D(n1731));   // src/ram.vhd(56[12:17])
    SB_DFF i2540_2541 (.Q(ram_s_105_2), .C(CLK_3P3_MHZ_c), .D(n1730));   // src/ram.vhd(56[12:17])
    SB_DFF i2537_2538 (.Q(ram_s_105_1), .C(CLK_3P3_MHZ_c), .D(n1729));   // src/ram.vhd(56[12:17])
    SB_DFF i2534_2535 (.Q(ram_s_105_0), .C(CLK_3P3_MHZ_c), .D(n1728));   // src/ram.vhd(56[12:17])
    SB_DFF i2531_2532 (.Q(ram_s_104_7), .C(CLK_3P3_MHZ_c), .D(n1727));   // src/ram.vhd(56[12:17])
    SB_DFF i2528_2529 (.Q(ram_s_104_6), .C(CLK_3P3_MHZ_c), .D(n1726));   // src/ram.vhd(56[12:17])
    SB_DFF i2525_2526 (.Q(ram_s_104_5), .C(CLK_3P3_MHZ_c), .D(n1725));   // src/ram.vhd(56[12:17])
    SB_DFF i2522_2523 (.Q(ram_s_104_4), .C(CLK_3P3_MHZ_c), .D(n1724));   // src/ram.vhd(56[12:17])
    SB_DFF i2519_2520 (.Q(ram_s_104_3), .C(CLK_3P3_MHZ_c), .D(n1723));   // src/ram.vhd(56[12:17])
    SB_DFF i2516_2517 (.Q(ram_s_104_2), .C(CLK_3P3_MHZ_c), .D(n1722));   // src/ram.vhd(56[12:17])
    SB_DFF i2513_2514 (.Q(ram_s_104_1), .C(CLK_3P3_MHZ_c), .D(n1721));   // src/ram.vhd(56[12:17])
    SB_DFF i2510_2511 (.Q(ram_s_104_0), .C(CLK_3P3_MHZ_c), .D(n1720));   // src/ram.vhd(56[12:17])
    SB_DFF i2507_2508 (.Q(ram_s_103_7), .C(CLK_3P3_MHZ_c), .D(n1719));   // src/ram.vhd(56[12:17])
    SB_DFF i2504_2505 (.Q(ram_s_103_6), .C(CLK_3P3_MHZ_c), .D(n1718));   // src/ram.vhd(56[12:17])
    SB_DFF i2501_2502 (.Q(ram_s_103_5), .C(CLK_3P3_MHZ_c), .D(n1717));   // src/ram.vhd(56[12:17])
    SB_DFF i2498_2499 (.Q(ram_s_103_4), .C(CLK_3P3_MHZ_c), .D(n1716));   // src/ram.vhd(56[12:17])
    SB_DFF i2495_2496 (.Q(ram_s_103_3), .C(CLK_3P3_MHZ_c), .D(n1715));   // src/ram.vhd(56[12:17])
    SB_DFF i2492_2493 (.Q(ram_s_103_2), .C(CLK_3P3_MHZ_c), .D(n1714));   // src/ram.vhd(56[12:17])
    SB_DFF i2489_2490 (.Q(ram_s_103_1), .C(CLK_3P3_MHZ_c), .D(n1713));   // src/ram.vhd(56[12:17])
    SB_DFF i2486_2487 (.Q(ram_s_103_0), .C(CLK_3P3_MHZ_c), .D(n1712));   // src/ram.vhd(56[12:17])
    SB_DFF i2483_2484 (.Q(ram_s_102_7), .C(CLK_3P3_MHZ_c), .D(n1711));   // src/ram.vhd(56[12:17])
    SB_DFF i2480_2481 (.Q(ram_s_102_6), .C(CLK_3P3_MHZ_c), .D(n1710));   // src/ram.vhd(56[12:17])
    SB_DFF i2477_2478 (.Q(ram_s_102_5), .C(CLK_3P3_MHZ_c), .D(n1709));   // src/ram.vhd(56[12:17])
    SB_DFF i2474_2475 (.Q(ram_s_102_4), .C(CLK_3P3_MHZ_c), .D(n1708));   // src/ram.vhd(56[12:17])
    SB_DFF i2471_2472 (.Q(ram_s_102_3), .C(CLK_3P3_MHZ_c), .D(n1707));   // src/ram.vhd(56[12:17])
    SB_DFF i2468_2469 (.Q(ram_s_102_2), .C(CLK_3P3_MHZ_c), .D(n1706));   // src/ram.vhd(56[12:17])
    SB_DFF i2465_2466 (.Q(ram_s_102_1), .C(CLK_3P3_MHZ_c), .D(n1705));   // src/ram.vhd(56[12:17])
    SB_DFF i2462_2463 (.Q(ram_s_102_0), .C(CLK_3P3_MHZ_c), .D(n1704));   // src/ram.vhd(56[12:17])
    SB_DFF i2459_2460 (.Q(ram_s_101_7), .C(CLK_3P3_MHZ_c), .D(n1703));   // src/ram.vhd(56[12:17])
    SB_DFF i2456_2457 (.Q(ram_s_101_6), .C(CLK_3P3_MHZ_c), .D(n1702));   // src/ram.vhd(56[12:17])
    SB_DFF i2453_2454 (.Q(ram_s_101_5), .C(CLK_3P3_MHZ_c), .D(n1701));   // src/ram.vhd(56[12:17])
    SB_DFF i2450_2451 (.Q(ram_s_101_4), .C(CLK_3P3_MHZ_c), .D(n1700));   // src/ram.vhd(56[12:17])
    SB_DFF i2447_2448 (.Q(ram_s_101_3), .C(CLK_3P3_MHZ_c), .D(n1699));   // src/ram.vhd(56[12:17])
    SB_DFF i2444_2445 (.Q(ram_s_101_2), .C(CLK_3P3_MHZ_c), .D(n1698));   // src/ram.vhd(56[12:17])
    SB_DFF i2441_2442 (.Q(ram_s_101_1), .C(CLK_3P3_MHZ_c), .D(n1697));   // src/ram.vhd(56[12:17])
    SB_DFF i2438_2439 (.Q(ram_s_101_0), .C(CLK_3P3_MHZ_c), .D(n1696));   // src/ram.vhd(56[12:17])
    SB_DFF i2435_2436 (.Q(ram_s_100_7), .C(CLK_3P3_MHZ_c), .D(n1695));   // src/ram.vhd(56[12:17])
    SB_DFF i2432_2433 (.Q(ram_s_100_6), .C(CLK_3P3_MHZ_c), .D(n1694));   // src/ram.vhd(56[12:17])
    SB_DFF i2429_2430 (.Q(ram_s_100_5), .C(CLK_3P3_MHZ_c), .D(n1693));   // src/ram.vhd(56[12:17])
    SB_DFF i2426_2427 (.Q(ram_s_100_4), .C(CLK_3P3_MHZ_c), .D(n1692));   // src/ram.vhd(56[12:17])
    SB_DFF i2423_2424 (.Q(ram_s_100_3), .C(CLK_3P3_MHZ_c), .D(n1691));   // src/ram.vhd(56[12:17])
    SB_DFF i2420_2421 (.Q(ram_s_100_2), .C(CLK_3P3_MHZ_c), .D(n1690));   // src/ram.vhd(56[12:17])
    SB_DFF i2417_2418 (.Q(ram_s_100_1), .C(CLK_3P3_MHZ_c), .D(n1689));   // src/ram.vhd(56[12:17])
    SB_DFF i2414_2415 (.Q(ram_s_100_0), .C(CLK_3P3_MHZ_c), .D(n1688));   // src/ram.vhd(56[12:17])
    SB_DFF i2411_2412 (.Q(ram_s_99_7), .C(CLK_3P3_MHZ_c), .D(n1687));   // src/ram.vhd(56[12:17])
    SB_DFF i2408_2409 (.Q(ram_s_99_6), .C(CLK_3P3_MHZ_c), .D(n1686));   // src/ram.vhd(56[12:17])
    SB_DFF i2405_2406 (.Q(ram_s_99_5), .C(CLK_3P3_MHZ_c), .D(n1685));   // src/ram.vhd(56[12:17])
    SB_DFF i2402_2403 (.Q(ram_s_99_4), .C(CLK_3P3_MHZ_c), .D(n1684));   // src/ram.vhd(56[12:17])
    SB_DFF i2399_2400 (.Q(ram_s_99_3), .C(CLK_3P3_MHZ_c), .D(n1683));   // src/ram.vhd(56[12:17])
    SB_DFF i2396_2397 (.Q(ram_s_99_2), .C(CLK_3P3_MHZ_c), .D(n1682));   // src/ram.vhd(56[12:17])
    SB_DFF i2393_2394 (.Q(ram_s_99_1), .C(CLK_3P3_MHZ_c), .D(n1681));   // src/ram.vhd(56[12:17])
    SB_DFF i2390_2391 (.Q(ram_s_99_0), .C(CLK_3P3_MHZ_c), .D(n1680));   // src/ram.vhd(56[12:17])
    SB_DFF i2387_2388 (.Q(ram_s_98_7), .C(CLK_3P3_MHZ_c), .D(n1679));   // src/ram.vhd(56[12:17])
    SB_DFF i2384_2385 (.Q(ram_s_98_6), .C(CLK_3P3_MHZ_c), .D(n1678));   // src/ram.vhd(56[12:17])
    SB_DFF i2381_2382 (.Q(ram_s_98_5), .C(CLK_3P3_MHZ_c), .D(n1677));   // src/ram.vhd(56[12:17])
    SB_DFF i2378_2379 (.Q(ram_s_98_4), .C(CLK_3P3_MHZ_c), .D(n1676));   // src/ram.vhd(56[12:17])
    SB_DFF i2375_2376 (.Q(ram_s_98_3), .C(CLK_3P3_MHZ_c), .D(n1675));   // src/ram.vhd(56[12:17])
    SB_DFF i2372_2373 (.Q(ram_s_98_2), .C(CLK_3P3_MHZ_c), .D(n1674));   // src/ram.vhd(56[12:17])
    SB_DFF i2369_2370 (.Q(ram_s_98_1), .C(CLK_3P3_MHZ_c), .D(n1673));   // src/ram.vhd(56[12:17])
    SB_DFF i2366_2367 (.Q(ram_s_98_0), .C(CLK_3P3_MHZ_c), .D(n1672));   // src/ram.vhd(56[12:17])
    SB_DFF i2363_2364 (.Q(ram_s_97_7), .C(CLK_3P3_MHZ_c), .D(n1671));   // src/ram.vhd(56[12:17])
    SB_DFF i2360_2361 (.Q(ram_s_97_6), .C(CLK_3P3_MHZ_c), .D(n1670));   // src/ram.vhd(56[12:17])
    SB_DFF i2357_2358 (.Q(ram_s_97_5), .C(CLK_3P3_MHZ_c), .D(n1669));   // src/ram.vhd(56[12:17])
    SB_DFF i2354_2355 (.Q(ram_s_97_4), .C(CLK_3P3_MHZ_c), .D(n1668));   // src/ram.vhd(56[12:17])
    SB_DFF i2351_2352 (.Q(ram_s_97_3), .C(CLK_3P3_MHZ_c), .D(n1667));   // src/ram.vhd(56[12:17])
    SB_DFF i2348_2349 (.Q(ram_s_97_2), .C(CLK_3P3_MHZ_c), .D(n1666));   // src/ram.vhd(56[12:17])
    SB_DFF i2345_2346 (.Q(ram_s_97_1), .C(CLK_3P3_MHZ_c), .D(n1665));   // src/ram.vhd(56[12:17])
    SB_DFF i2342_2343 (.Q(ram_s_97_0), .C(CLK_3P3_MHZ_c), .D(n1664));   // src/ram.vhd(56[12:17])
    SB_DFF i2339_2340 (.Q(ram_s_96_7), .C(CLK_3P3_MHZ_c), .D(n1663));   // src/ram.vhd(56[12:17])
    SB_DFF i2336_2337 (.Q(ram_s_96_6), .C(CLK_3P3_MHZ_c), .D(n1662));   // src/ram.vhd(56[12:17])
    SB_DFF i2333_2334 (.Q(ram_s_96_5), .C(CLK_3P3_MHZ_c), .D(n1661));   // src/ram.vhd(56[12:17])
    SB_DFF i2330_2331 (.Q(ram_s_96_4), .C(CLK_3P3_MHZ_c), .D(n1660));   // src/ram.vhd(56[12:17])
    SB_DFF i2327_2328 (.Q(ram_s_96_3), .C(CLK_3P3_MHZ_c), .D(n1659));   // src/ram.vhd(56[12:17])
    SB_DFF i2324_2325 (.Q(ram_s_96_2), .C(CLK_3P3_MHZ_c), .D(n1658));   // src/ram.vhd(56[12:17])
    SB_DFF i2321_2322 (.Q(ram_s_96_1), .C(CLK_3P3_MHZ_c), .D(n1657));   // src/ram.vhd(56[12:17])
    SB_DFF i2318_2319 (.Q(ram_s_96_0), .C(CLK_3P3_MHZ_c), .D(n1656));   // src/ram.vhd(56[12:17])
    SB_DFF i2315_2316 (.Q(ram_s_95_7), .C(CLK_3P3_MHZ_c), .D(n1655));   // src/ram.vhd(56[12:17])
    SB_DFF i2312_2313 (.Q(ram_s_95_6), .C(CLK_3P3_MHZ_c), .D(n1654));   // src/ram.vhd(56[12:17])
    SB_DFF i2309_2310 (.Q(ram_s_95_5), .C(CLK_3P3_MHZ_c), .D(n1653));   // src/ram.vhd(56[12:17])
    SB_DFF i2306_2307 (.Q(ram_s_95_4), .C(CLK_3P3_MHZ_c), .D(n1652));   // src/ram.vhd(56[12:17])
    SB_DFF i2303_2304 (.Q(ram_s_95_3), .C(CLK_3P3_MHZ_c), .D(n1651));   // src/ram.vhd(56[12:17])
    SB_DFF i2300_2301 (.Q(ram_s_95_2), .C(CLK_3P3_MHZ_c), .D(n1650));   // src/ram.vhd(56[12:17])
    SB_DFF i2297_2298 (.Q(ram_s_95_1), .C(CLK_3P3_MHZ_c), .D(n1649));   // src/ram.vhd(56[12:17])
    SB_DFF i2294_2295 (.Q(ram_s_95_0), .C(CLK_3P3_MHZ_c), .D(n1648));   // src/ram.vhd(56[12:17])
    SB_DFF i2291_2292 (.Q(ram_s_94_7), .C(CLK_3P3_MHZ_c), .D(n1647));   // src/ram.vhd(56[12:17])
    SB_DFF i2288_2289 (.Q(ram_s_94_6), .C(CLK_3P3_MHZ_c), .D(n1646));   // src/ram.vhd(56[12:17])
    SB_DFF i2285_2286 (.Q(ram_s_94_5), .C(CLK_3P3_MHZ_c), .D(n1645));   // src/ram.vhd(56[12:17])
    SB_DFF i2282_2283 (.Q(ram_s_94_4), .C(CLK_3P3_MHZ_c), .D(n1644));   // src/ram.vhd(56[12:17])
    SB_DFF i2279_2280 (.Q(ram_s_94_3), .C(CLK_3P3_MHZ_c), .D(n1643));   // src/ram.vhd(56[12:17])
    SB_DFF i2276_2277 (.Q(ram_s_94_2), .C(CLK_3P3_MHZ_c), .D(n1642));   // src/ram.vhd(56[12:17])
    SB_DFF i2273_2274 (.Q(ram_s_94_1), .C(CLK_3P3_MHZ_c), .D(n1641));   // src/ram.vhd(56[12:17])
    SB_DFF i2270_2271 (.Q(ram_s_94_0), .C(CLK_3P3_MHZ_c), .D(n1640));   // src/ram.vhd(56[12:17])
    SB_DFF i2267_2268 (.Q(ram_s_93_7), .C(CLK_3P3_MHZ_c), .D(n1639));   // src/ram.vhd(56[12:17])
    SB_DFF i2264_2265 (.Q(ram_s_93_6), .C(CLK_3P3_MHZ_c), .D(n1638));   // src/ram.vhd(56[12:17])
    SB_DFF i2261_2262 (.Q(ram_s_93_5), .C(CLK_3P3_MHZ_c), .D(n1637));   // src/ram.vhd(56[12:17])
    SB_DFF i2258_2259 (.Q(ram_s_93_4), .C(CLK_3P3_MHZ_c), .D(n1636));   // src/ram.vhd(56[12:17])
    SB_DFF i2255_2256 (.Q(ram_s_93_3), .C(CLK_3P3_MHZ_c), .D(n1635));   // src/ram.vhd(56[12:17])
    SB_DFF i2252_2253 (.Q(ram_s_93_2), .C(CLK_3P3_MHZ_c), .D(n1634));   // src/ram.vhd(56[12:17])
    SB_DFF i2249_2250 (.Q(ram_s_93_1), .C(CLK_3P3_MHZ_c), .D(n1633));   // src/ram.vhd(56[12:17])
    SB_DFF i2246_2247 (.Q(ram_s_93_0), .C(CLK_3P3_MHZ_c), .D(n1632));   // src/ram.vhd(56[12:17])
    SB_DFF i2243_2244 (.Q(ram_s_92_7), .C(CLK_3P3_MHZ_c), .D(n1631));   // src/ram.vhd(56[12:17])
    SB_DFF i2240_2241 (.Q(ram_s_92_6), .C(CLK_3P3_MHZ_c), .D(n1630));   // src/ram.vhd(56[12:17])
    SB_DFF i2237_2238 (.Q(ram_s_92_5), .C(CLK_3P3_MHZ_c), .D(n1629));   // src/ram.vhd(56[12:17])
    SB_DFF i2234_2235 (.Q(ram_s_92_4), .C(CLK_3P3_MHZ_c), .D(n1628));   // src/ram.vhd(56[12:17])
    SB_DFF i2231_2232 (.Q(ram_s_92_3), .C(CLK_3P3_MHZ_c), .D(n1627));   // src/ram.vhd(56[12:17])
    SB_DFF i2228_2229 (.Q(ram_s_92_2), .C(CLK_3P3_MHZ_c), .D(n1626));   // src/ram.vhd(56[12:17])
    SB_DFF i2225_2226 (.Q(ram_s_92_1), .C(CLK_3P3_MHZ_c), .D(n1625));   // src/ram.vhd(56[12:17])
    SB_DFF i2222_2223 (.Q(ram_s_92_0), .C(CLK_3P3_MHZ_c), .D(n1624));   // src/ram.vhd(56[12:17])
    SB_DFF i2219_2220 (.Q(ram_s_91_7), .C(CLK_3P3_MHZ_c), .D(n1623));   // src/ram.vhd(56[12:17])
    SB_DFF i2216_2217 (.Q(ram_s_91_6), .C(CLK_3P3_MHZ_c), .D(n1622));   // src/ram.vhd(56[12:17])
    SB_DFF i2213_2214 (.Q(ram_s_91_5), .C(CLK_3P3_MHZ_c), .D(n1621));   // src/ram.vhd(56[12:17])
    SB_DFF i2210_2211 (.Q(ram_s_91_4), .C(CLK_3P3_MHZ_c), .D(n1620));   // src/ram.vhd(56[12:17])
    SB_DFF i2207_2208 (.Q(ram_s_91_3), .C(CLK_3P3_MHZ_c), .D(n1619));   // src/ram.vhd(56[12:17])
    SB_DFF i2204_2205 (.Q(ram_s_91_2), .C(CLK_3P3_MHZ_c), .D(n1618));   // src/ram.vhd(56[12:17])
    SB_DFF i2201_2202 (.Q(ram_s_91_1), .C(CLK_3P3_MHZ_c), .D(n1617));   // src/ram.vhd(56[12:17])
    SB_DFF i2198_2199 (.Q(ram_s_91_0), .C(CLK_3P3_MHZ_c), .D(n1616));   // src/ram.vhd(56[12:17])
    SB_DFF i2195_2196 (.Q(ram_s_90_7), .C(CLK_3P3_MHZ_c), .D(n1615));   // src/ram.vhd(56[12:17])
    SB_DFF i2192_2193 (.Q(ram_s_90_6), .C(CLK_3P3_MHZ_c), .D(n1614));   // src/ram.vhd(56[12:17])
    SB_DFF i2189_2190 (.Q(ram_s_90_5), .C(CLK_3P3_MHZ_c), .D(n1613));   // src/ram.vhd(56[12:17])
    SB_DFF i2186_2187 (.Q(ram_s_90_4), .C(CLK_3P3_MHZ_c), .D(n1612));   // src/ram.vhd(56[12:17])
    SB_DFF i2183_2184 (.Q(ram_s_90_3), .C(CLK_3P3_MHZ_c), .D(n1611));   // src/ram.vhd(56[12:17])
    SB_DFF i2180_2181 (.Q(ram_s_90_2), .C(CLK_3P3_MHZ_c), .D(n1610));   // src/ram.vhd(56[12:17])
    SB_DFF i2177_2178 (.Q(ram_s_90_1), .C(CLK_3P3_MHZ_c), .D(n1609));   // src/ram.vhd(56[12:17])
    SB_DFF i2174_2175 (.Q(ram_s_90_0), .C(CLK_3P3_MHZ_c), .D(n1608));   // src/ram.vhd(56[12:17])
    SB_DFF i2171_2172 (.Q(ram_s_89_7), .C(CLK_3P3_MHZ_c), .D(n1607));   // src/ram.vhd(56[12:17])
    SB_DFF i2168_2169 (.Q(ram_s_89_6), .C(CLK_3P3_MHZ_c), .D(n1606));   // src/ram.vhd(56[12:17])
    SB_DFF i2165_2166 (.Q(ram_s_89_5), .C(CLK_3P3_MHZ_c), .D(n1605));   // src/ram.vhd(56[12:17])
    SB_DFF i2162_2163 (.Q(ram_s_89_4), .C(CLK_3P3_MHZ_c), .D(n1604));   // src/ram.vhd(56[12:17])
    SB_DFF i2159_2160 (.Q(ram_s_89_3), .C(CLK_3P3_MHZ_c), .D(n1603));   // src/ram.vhd(56[12:17])
    SB_DFF i2156_2157 (.Q(ram_s_89_2), .C(CLK_3P3_MHZ_c), .D(n1602));   // src/ram.vhd(56[12:17])
    SB_DFF i2153_2154 (.Q(ram_s_89_1), .C(CLK_3P3_MHZ_c), .D(n1601));   // src/ram.vhd(56[12:17])
    SB_DFF i2150_2151 (.Q(ram_s_89_0), .C(CLK_3P3_MHZ_c), .D(n1600));   // src/ram.vhd(56[12:17])
    SB_DFF i2147_2148 (.Q(ram_s_88_7), .C(CLK_3P3_MHZ_c), .D(n1599));   // src/ram.vhd(56[12:17])
    SB_DFF i2144_2145 (.Q(ram_s_88_6), .C(CLK_3P3_MHZ_c), .D(n1598));   // src/ram.vhd(56[12:17])
    SB_DFF i2141_2142 (.Q(ram_s_88_5), .C(CLK_3P3_MHZ_c), .D(n1597));   // src/ram.vhd(56[12:17])
    SB_DFF i2138_2139 (.Q(ram_s_88_4), .C(CLK_3P3_MHZ_c), .D(n1596));   // src/ram.vhd(56[12:17])
    SB_DFF i2135_2136 (.Q(ram_s_88_3), .C(CLK_3P3_MHZ_c), .D(n1595));   // src/ram.vhd(56[12:17])
    SB_DFF i2132_2133 (.Q(ram_s_88_2), .C(CLK_3P3_MHZ_c), .D(n1594));   // src/ram.vhd(56[12:17])
    SB_DFF i2129_2130 (.Q(ram_s_88_1), .C(CLK_3P3_MHZ_c), .D(n1593));   // src/ram.vhd(56[12:17])
    SB_DFF i2126_2127 (.Q(ram_s_88_0), .C(CLK_3P3_MHZ_c), .D(n1592));   // src/ram.vhd(56[12:17])
    SB_DFF i2123_2124 (.Q(ram_s_87_7), .C(CLK_3P3_MHZ_c), .D(n1591));   // src/ram.vhd(56[12:17])
    SB_DFF i2120_2121 (.Q(ram_s_87_6), .C(CLK_3P3_MHZ_c), .D(n1590));   // src/ram.vhd(56[12:17])
    SB_DFF i2117_2118 (.Q(ram_s_87_5), .C(CLK_3P3_MHZ_c), .D(n1589));   // src/ram.vhd(56[12:17])
    SB_DFF i2114_2115 (.Q(ram_s_87_4), .C(CLK_3P3_MHZ_c), .D(n1588));   // src/ram.vhd(56[12:17])
    SB_DFF i2111_2112 (.Q(ram_s_87_3), .C(CLK_3P3_MHZ_c), .D(n1587));   // src/ram.vhd(56[12:17])
    SB_DFF i2108_2109 (.Q(ram_s_87_2), .C(CLK_3P3_MHZ_c), .D(n1586));   // src/ram.vhd(56[12:17])
    SB_DFF i2105_2106 (.Q(ram_s_87_1), .C(CLK_3P3_MHZ_c), .D(n1585));   // src/ram.vhd(56[12:17])
    SB_DFF i2102_2103 (.Q(ram_s_87_0), .C(CLK_3P3_MHZ_c), .D(n1584));   // src/ram.vhd(56[12:17])
    SB_DFF i2099_2100 (.Q(ram_s_86_7), .C(CLK_3P3_MHZ_c), .D(n1583));   // src/ram.vhd(56[12:17])
    SB_DFF i2096_2097 (.Q(ram_s_86_6), .C(CLK_3P3_MHZ_c), .D(n1582));   // src/ram.vhd(56[12:17])
    SB_DFF i2093_2094 (.Q(ram_s_86_5), .C(CLK_3P3_MHZ_c), .D(n1581));   // src/ram.vhd(56[12:17])
    SB_DFF i2090_2091 (.Q(ram_s_86_4), .C(CLK_3P3_MHZ_c), .D(n1580));   // src/ram.vhd(56[12:17])
    SB_DFF i2087_2088 (.Q(ram_s_86_3), .C(CLK_3P3_MHZ_c), .D(n1579));   // src/ram.vhd(56[12:17])
    SB_DFF i2084_2085 (.Q(ram_s_86_2), .C(CLK_3P3_MHZ_c), .D(n1578));   // src/ram.vhd(56[12:17])
    SB_DFF i2081_2082 (.Q(ram_s_86_1), .C(CLK_3P3_MHZ_c), .D(n1577));   // src/ram.vhd(56[12:17])
    SB_DFF i2078_2079 (.Q(ram_s_86_0), .C(CLK_3P3_MHZ_c), .D(n1576));   // src/ram.vhd(56[12:17])
    SB_DFF i2075_2076 (.Q(ram_s_85_7), .C(CLK_3P3_MHZ_c), .D(n1575));   // src/ram.vhd(56[12:17])
    SB_DFF i2072_2073 (.Q(ram_s_85_6), .C(CLK_3P3_MHZ_c), .D(n1574));   // src/ram.vhd(56[12:17])
    SB_DFF i2069_2070 (.Q(ram_s_85_5), .C(CLK_3P3_MHZ_c), .D(n1573));   // src/ram.vhd(56[12:17])
    SB_DFF i2066_2067 (.Q(ram_s_85_4), .C(CLK_3P3_MHZ_c), .D(n1572));   // src/ram.vhd(56[12:17])
    SB_DFF i2063_2064 (.Q(ram_s_85_3), .C(CLK_3P3_MHZ_c), .D(n1571));   // src/ram.vhd(56[12:17])
    SB_DFF i2060_2061 (.Q(ram_s_85_2), .C(CLK_3P3_MHZ_c), .D(n1570));   // src/ram.vhd(56[12:17])
    SB_DFF i2057_2058 (.Q(ram_s_85_1), .C(CLK_3P3_MHZ_c), .D(n1569));   // src/ram.vhd(56[12:17])
    SB_DFF i2054_2055 (.Q(ram_s_85_0), .C(CLK_3P3_MHZ_c), .D(n1568));   // src/ram.vhd(56[12:17])
    SB_DFF i2051_2052 (.Q(ram_s_84_7), .C(CLK_3P3_MHZ_c), .D(n1567));   // src/ram.vhd(56[12:17])
    SB_DFF i2048_2049 (.Q(ram_s_84_6), .C(CLK_3P3_MHZ_c), .D(n1566));   // src/ram.vhd(56[12:17])
    SB_DFF i2045_2046 (.Q(ram_s_84_5), .C(CLK_3P3_MHZ_c), .D(n1565));   // src/ram.vhd(56[12:17])
    SB_DFF i2042_2043 (.Q(ram_s_84_4), .C(CLK_3P3_MHZ_c), .D(n1564));   // src/ram.vhd(56[12:17])
    SB_DFF i2039_2040 (.Q(ram_s_84_3), .C(CLK_3P3_MHZ_c), .D(n1563));   // src/ram.vhd(56[12:17])
    SB_DFF i2036_2037 (.Q(ram_s_84_2), .C(CLK_3P3_MHZ_c), .D(n1562));   // src/ram.vhd(56[12:17])
    SB_DFF i2033_2034 (.Q(ram_s_84_1), .C(CLK_3P3_MHZ_c), .D(n1561));   // src/ram.vhd(56[12:17])
    SB_DFF i2030_2031 (.Q(ram_s_84_0), .C(CLK_3P3_MHZ_c), .D(n1560));   // src/ram.vhd(56[12:17])
    SB_DFF i2027_2028 (.Q(ram_s_83_7), .C(CLK_3P3_MHZ_c), .D(n1559));   // src/ram.vhd(56[12:17])
    SB_DFF i2024_2025 (.Q(ram_s_83_6), .C(CLK_3P3_MHZ_c), .D(n1558));   // src/ram.vhd(56[12:17])
    SB_DFF i2021_2022 (.Q(ram_s_83_5), .C(CLK_3P3_MHZ_c), .D(n1557));   // src/ram.vhd(56[12:17])
    SB_DFF i2018_2019 (.Q(ram_s_83_4), .C(CLK_3P3_MHZ_c), .D(n1556));   // src/ram.vhd(56[12:17])
    SB_DFF i2015_2016 (.Q(ram_s_83_3), .C(CLK_3P3_MHZ_c), .D(n1555));   // src/ram.vhd(56[12:17])
    SB_DFF i2012_2013 (.Q(ram_s_83_2), .C(CLK_3P3_MHZ_c), .D(n1554));   // src/ram.vhd(56[12:17])
    SB_DFF i2009_2010 (.Q(ram_s_83_1), .C(CLK_3P3_MHZ_c), .D(n1553));   // src/ram.vhd(56[12:17])
    SB_DFF i2006_2007 (.Q(ram_s_83_0), .C(CLK_3P3_MHZ_c), .D(n1552));   // src/ram.vhd(56[12:17])
    SB_DFF i2003_2004 (.Q(ram_s_82_7), .C(CLK_3P3_MHZ_c), .D(n1551));   // src/ram.vhd(56[12:17])
    SB_DFF i2000_2001 (.Q(ram_s_82_6), .C(CLK_3P3_MHZ_c), .D(n1550));   // src/ram.vhd(56[12:17])
    SB_DFF i1997_1998 (.Q(ram_s_82_5), .C(CLK_3P3_MHZ_c), .D(n1549));   // src/ram.vhd(56[12:17])
    SB_DFF i1994_1995 (.Q(ram_s_82_4), .C(CLK_3P3_MHZ_c), .D(n1548));   // src/ram.vhd(56[12:17])
    SB_DFF i1991_1992 (.Q(ram_s_82_3), .C(CLK_3P3_MHZ_c), .D(n1547));   // src/ram.vhd(56[12:17])
    SB_DFF i1988_1989 (.Q(ram_s_82_2), .C(CLK_3P3_MHZ_c), .D(n1546));   // src/ram.vhd(56[12:17])
    SB_DFF i1985_1986 (.Q(ram_s_82_1), .C(CLK_3P3_MHZ_c), .D(n1545));   // src/ram.vhd(56[12:17])
    SB_DFF i1982_1983 (.Q(ram_s_82_0), .C(CLK_3P3_MHZ_c), .D(n1544));   // src/ram.vhd(56[12:17])
    SB_DFF i1979_1980 (.Q(ram_s_81_7), .C(CLK_3P3_MHZ_c), .D(n1543));   // src/ram.vhd(56[12:17])
    SB_DFF i1976_1977 (.Q(ram_s_81_6), .C(CLK_3P3_MHZ_c), .D(n1542));   // src/ram.vhd(56[12:17])
    SB_DFF i1973_1974 (.Q(ram_s_81_5), .C(CLK_3P3_MHZ_c), .D(n1541));   // src/ram.vhd(56[12:17])
    SB_DFF i1970_1971 (.Q(ram_s_81_4), .C(CLK_3P3_MHZ_c), .D(n1540));   // src/ram.vhd(56[12:17])
    SB_DFF i1967_1968 (.Q(ram_s_81_3), .C(CLK_3P3_MHZ_c), .D(n1539));   // src/ram.vhd(56[12:17])
    SB_DFF i1964_1965 (.Q(ram_s_81_2), .C(CLK_3P3_MHZ_c), .D(n1538));   // src/ram.vhd(56[12:17])
    SB_DFF i1961_1962 (.Q(ram_s_81_1), .C(CLK_3P3_MHZ_c), .D(n1537));   // src/ram.vhd(56[12:17])
    SB_DFF i1958_1959 (.Q(ram_s_81_0), .C(CLK_3P3_MHZ_c), .D(n1536));   // src/ram.vhd(56[12:17])
    SB_DFF i1955_1956 (.Q(ram_s_80_7), .C(CLK_3P3_MHZ_c), .D(n1535));   // src/ram.vhd(56[12:17])
    SB_DFF i1952_1953 (.Q(ram_s_80_6), .C(CLK_3P3_MHZ_c), .D(n1534));   // src/ram.vhd(56[12:17])
    SB_DFF i1949_1950 (.Q(ram_s_80_5), .C(CLK_3P3_MHZ_c), .D(n1533));   // src/ram.vhd(56[12:17])
    SB_DFF i1946_1947 (.Q(ram_s_80_4), .C(CLK_3P3_MHZ_c), .D(n1532));   // src/ram.vhd(56[12:17])
    SB_DFF i1943_1944 (.Q(ram_s_80_3), .C(CLK_3P3_MHZ_c), .D(n1531));   // src/ram.vhd(56[12:17])
    SB_DFF i1940_1941 (.Q(ram_s_80_2), .C(CLK_3P3_MHZ_c), .D(n1530));   // src/ram.vhd(56[12:17])
    SB_DFF i1937_1938 (.Q(ram_s_80_1), .C(CLK_3P3_MHZ_c), .D(n1529));   // src/ram.vhd(56[12:17])
    SB_DFF i1934_1935 (.Q(ram_s_80_0), .C(CLK_3P3_MHZ_c), .D(n1528));   // src/ram.vhd(56[12:17])
    SB_DFF i1931_1932 (.Q(ram_s_79_7), .C(CLK_3P3_MHZ_c), .D(n1527));   // src/ram.vhd(56[12:17])
    SB_DFF i1928_1929 (.Q(ram_s_79_6), .C(CLK_3P3_MHZ_c), .D(n1526));   // src/ram.vhd(56[12:17])
    SB_DFF i1925_1926 (.Q(ram_s_79_5), .C(CLK_3P3_MHZ_c), .D(n1525));   // src/ram.vhd(56[12:17])
    SB_DFF i1922_1923 (.Q(ram_s_79_4), .C(CLK_3P3_MHZ_c), .D(n1524));   // src/ram.vhd(56[12:17])
    SB_DFF i1919_1920 (.Q(ram_s_79_3), .C(CLK_3P3_MHZ_c), .D(n1523));   // src/ram.vhd(56[12:17])
    SB_DFF i1916_1917 (.Q(ram_s_79_2), .C(CLK_3P3_MHZ_c), .D(n1522));   // src/ram.vhd(56[12:17])
    SB_DFF i1913_1914 (.Q(ram_s_79_1), .C(CLK_3P3_MHZ_c), .D(n1521));   // src/ram.vhd(56[12:17])
    SB_DFF i1910_1911 (.Q(ram_s_79_0), .C(CLK_3P3_MHZ_c), .D(n1520));   // src/ram.vhd(56[12:17])
    SB_DFF i1907_1908 (.Q(ram_s_78_7), .C(CLK_3P3_MHZ_c), .D(n1519));   // src/ram.vhd(56[12:17])
    SB_DFF i1904_1905 (.Q(ram_s_78_6), .C(CLK_3P3_MHZ_c), .D(n1518));   // src/ram.vhd(56[12:17])
    SB_DFF i1901_1902 (.Q(ram_s_78_5), .C(CLK_3P3_MHZ_c), .D(n1517));   // src/ram.vhd(56[12:17])
    SB_DFF i1898_1899 (.Q(ram_s_78_4), .C(CLK_3P3_MHZ_c), .D(n1516));   // src/ram.vhd(56[12:17])
    SB_DFF i1895_1896 (.Q(ram_s_78_3), .C(CLK_3P3_MHZ_c), .D(n1515));   // src/ram.vhd(56[12:17])
    SB_DFF i1892_1893 (.Q(ram_s_78_2), .C(CLK_3P3_MHZ_c), .D(n1514));   // src/ram.vhd(56[12:17])
    SB_DFF i1889_1890 (.Q(ram_s_78_1), .C(CLK_3P3_MHZ_c), .D(n1513));   // src/ram.vhd(56[12:17])
    SB_DFF i1886_1887 (.Q(ram_s_78_0), .C(CLK_3P3_MHZ_c), .D(n1512));   // src/ram.vhd(56[12:17])
    SB_DFF i1883_1884 (.Q(ram_s_77_7), .C(CLK_3P3_MHZ_c), .D(n1511));   // src/ram.vhd(56[12:17])
    SB_DFF i1880_1881 (.Q(ram_s_77_6), .C(CLK_3P3_MHZ_c), .D(n1510));   // src/ram.vhd(56[12:17])
    SB_DFF i1877_1878 (.Q(ram_s_77_5), .C(CLK_3P3_MHZ_c), .D(n1509));   // src/ram.vhd(56[12:17])
    SB_DFF i1874_1875 (.Q(ram_s_77_4), .C(CLK_3P3_MHZ_c), .D(n1508));   // src/ram.vhd(56[12:17])
    SB_DFF i1871_1872 (.Q(ram_s_77_3), .C(CLK_3P3_MHZ_c), .D(n1507));   // src/ram.vhd(56[12:17])
    SB_DFF i1868_1869 (.Q(ram_s_77_2), .C(CLK_3P3_MHZ_c), .D(n1506));   // src/ram.vhd(56[12:17])
    SB_DFF i1865_1866 (.Q(ram_s_77_1), .C(CLK_3P3_MHZ_c), .D(n1505));   // src/ram.vhd(56[12:17])
    SB_DFF i1862_1863 (.Q(ram_s_77_0), .C(CLK_3P3_MHZ_c), .D(n1504));   // src/ram.vhd(56[12:17])
    SB_DFF i1859_1860 (.Q(ram_s_76_7), .C(CLK_3P3_MHZ_c), .D(n1503));   // src/ram.vhd(56[12:17])
    SB_DFF i1856_1857 (.Q(ram_s_76_6), .C(CLK_3P3_MHZ_c), .D(n1502));   // src/ram.vhd(56[12:17])
    SB_DFF i1853_1854 (.Q(ram_s_76_5), .C(CLK_3P3_MHZ_c), .D(n1501));   // src/ram.vhd(56[12:17])
    SB_DFF i1850_1851 (.Q(ram_s_76_4), .C(CLK_3P3_MHZ_c), .D(n1500));   // src/ram.vhd(56[12:17])
    SB_DFF i1847_1848 (.Q(ram_s_76_3), .C(CLK_3P3_MHZ_c), .D(n1499));   // src/ram.vhd(56[12:17])
    SB_DFF i1844_1845 (.Q(ram_s_76_2), .C(CLK_3P3_MHZ_c), .D(n1498));   // src/ram.vhd(56[12:17])
    SB_DFF i1841_1842 (.Q(ram_s_76_1), .C(CLK_3P3_MHZ_c), .D(n1497));   // src/ram.vhd(56[12:17])
    SB_DFF i1838_1839 (.Q(ram_s_76_0), .C(CLK_3P3_MHZ_c), .D(n1496));   // src/ram.vhd(56[12:17])
    SB_DFF i1835_1836 (.Q(ram_s_75_7), .C(CLK_3P3_MHZ_c), .D(n1495));   // src/ram.vhd(56[12:17])
    SB_DFF i1832_1833 (.Q(ram_s_75_6), .C(CLK_3P3_MHZ_c), .D(n1494));   // src/ram.vhd(56[12:17])
    SB_DFF i1829_1830 (.Q(ram_s_75_5), .C(CLK_3P3_MHZ_c), .D(n1493));   // src/ram.vhd(56[12:17])
    SB_DFF i1826_1827 (.Q(ram_s_75_4), .C(CLK_3P3_MHZ_c), .D(n1492));   // src/ram.vhd(56[12:17])
    SB_DFF i1823_1824 (.Q(ram_s_75_3), .C(CLK_3P3_MHZ_c), .D(n1491));   // src/ram.vhd(56[12:17])
    SB_DFF i1820_1821 (.Q(ram_s_75_2), .C(CLK_3P3_MHZ_c), .D(n1490));   // src/ram.vhd(56[12:17])
    SB_DFF i1817_1818 (.Q(ram_s_75_1), .C(CLK_3P3_MHZ_c), .D(n1489));   // src/ram.vhd(56[12:17])
    SB_DFF i1814_1815 (.Q(ram_s_75_0), .C(CLK_3P3_MHZ_c), .D(n1488));   // src/ram.vhd(56[12:17])
    SB_DFF i1811_1812 (.Q(ram_s_74_7), .C(CLK_3P3_MHZ_c), .D(n1487));   // src/ram.vhd(56[12:17])
    SB_DFF i1808_1809 (.Q(ram_s_74_6), .C(CLK_3P3_MHZ_c), .D(n1486));   // src/ram.vhd(56[12:17])
    SB_DFF i1805_1806 (.Q(ram_s_74_5), .C(CLK_3P3_MHZ_c), .D(n1485));   // src/ram.vhd(56[12:17])
    SB_DFF i1802_1803 (.Q(ram_s_74_4), .C(CLK_3P3_MHZ_c), .D(n1484));   // src/ram.vhd(56[12:17])
    SB_DFF i1799_1800 (.Q(ram_s_74_3), .C(CLK_3P3_MHZ_c), .D(n1483));   // src/ram.vhd(56[12:17])
    SB_DFF i1796_1797 (.Q(ram_s_74_2), .C(CLK_3P3_MHZ_c), .D(n1482));   // src/ram.vhd(56[12:17])
    SB_DFF i1793_1794 (.Q(ram_s_74_1), .C(CLK_3P3_MHZ_c), .D(n1481));   // src/ram.vhd(56[12:17])
    SB_DFF i1790_1791 (.Q(ram_s_74_0), .C(CLK_3P3_MHZ_c), .D(n1480));   // src/ram.vhd(56[12:17])
    SB_DFF i1787_1788 (.Q(ram_s_73_7), .C(CLK_3P3_MHZ_c), .D(n1479));   // src/ram.vhd(56[12:17])
    SB_DFF i1784_1785 (.Q(ram_s_73_6), .C(CLK_3P3_MHZ_c), .D(n1478));   // src/ram.vhd(56[12:17])
    SB_DFF i1781_1782 (.Q(ram_s_73_5), .C(CLK_3P3_MHZ_c), .D(n1477));   // src/ram.vhd(56[12:17])
    SB_DFF i1778_1779 (.Q(ram_s_73_4), .C(CLK_3P3_MHZ_c), .D(n1476));   // src/ram.vhd(56[12:17])
    SB_DFF i1775_1776 (.Q(ram_s_73_3), .C(CLK_3P3_MHZ_c), .D(n1475));   // src/ram.vhd(56[12:17])
    SB_DFF i1772_1773 (.Q(ram_s_73_2), .C(CLK_3P3_MHZ_c), .D(n1474));   // src/ram.vhd(56[12:17])
    SB_DFF i1769_1770 (.Q(ram_s_73_1), .C(CLK_3P3_MHZ_c), .D(n1473));   // src/ram.vhd(56[12:17])
    SB_DFF i1766_1767 (.Q(ram_s_73_0), .C(CLK_3P3_MHZ_c), .D(n1472));   // src/ram.vhd(56[12:17])
    SB_DFF i1763_1764 (.Q(ram_s_72_7), .C(CLK_3P3_MHZ_c), .D(n1471));   // src/ram.vhd(56[12:17])
    SB_DFF i1760_1761 (.Q(ram_s_72_6), .C(CLK_3P3_MHZ_c), .D(n1470));   // src/ram.vhd(56[12:17])
    SB_DFF i1757_1758 (.Q(ram_s_72_5), .C(CLK_3P3_MHZ_c), .D(n1469));   // src/ram.vhd(56[12:17])
    SB_DFF i1754_1755 (.Q(ram_s_72_4), .C(CLK_3P3_MHZ_c), .D(n1468));   // src/ram.vhd(56[12:17])
    SB_DFF i1751_1752 (.Q(ram_s_72_3), .C(CLK_3P3_MHZ_c), .D(n1467));   // src/ram.vhd(56[12:17])
    SB_DFF i1748_1749 (.Q(ram_s_72_2), .C(CLK_3P3_MHZ_c), .D(n1466));   // src/ram.vhd(56[12:17])
    SB_DFF i1745_1746 (.Q(ram_s_72_1), .C(CLK_3P3_MHZ_c), .D(n1465));   // src/ram.vhd(56[12:17])
    SB_DFF i1742_1743 (.Q(ram_s_72_0), .C(CLK_3P3_MHZ_c), .D(n1464));   // src/ram.vhd(56[12:17])
    SB_DFF i1739_1740 (.Q(ram_s_71_7), .C(CLK_3P3_MHZ_c), .D(n1463));   // src/ram.vhd(56[12:17])
    SB_DFF i1736_1737 (.Q(ram_s_71_6), .C(CLK_3P3_MHZ_c), .D(n1462));   // src/ram.vhd(56[12:17])
    SB_DFF i1733_1734 (.Q(ram_s_71_5), .C(CLK_3P3_MHZ_c), .D(n1461));   // src/ram.vhd(56[12:17])
    SB_DFF i1730_1731 (.Q(ram_s_71_4), .C(CLK_3P3_MHZ_c), .D(n1460));   // src/ram.vhd(56[12:17])
    SB_DFF i1727_1728 (.Q(ram_s_71_3), .C(CLK_3P3_MHZ_c), .D(n1459));   // src/ram.vhd(56[12:17])
    SB_DFF i1724_1725 (.Q(ram_s_71_2), .C(CLK_3P3_MHZ_c), .D(n1458));   // src/ram.vhd(56[12:17])
    SB_DFF i1721_1722 (.Q(ram_s_71_1), .C(CLK_3P3_MHZ_c), .D(n1457));   // src/ram.vhd(56[12:17])
    SB_DFF i1718_1719 (.Q(ram_s_71_0), .C(CLK_3P3_MHZ_c), .D(n1456));   // src/ram.vhd(56[12:17])
    SB_DFF i1715_1716 (.Q(ram_s_70_7), .C(CLK_3P3_MHZ_c), .D(n1455));   // src/ram.vhd(56[12:17])
    SB_DFF i1712_1713 (.Q(ram_s_70_6), .C(CLK_3P3_MHZ_c), .D(n1454));   // src/ram.vhd(56[12:17])
    SB_DFF i1709_1710 (.Q(ram_s_70_5), .C(CLK_3P3_MHZ_c), .D(n1453));   // src/ram.vhd(56[12:17])
    SB_DFF i1706_1707 (.Q(ram_s_70_4), .C(CLK_3P3_MHZ_c), .D(n1452));   // src/ram.vhd(56[12:17])
    SB_DFF i1703_1704 (.Q(ram_s_70_3), .C(CLK_3P3_MHZ_c), .D(n1451));   // src/ram.vhd(56[12:17])
    SB_DFF i1700_1701 (.Q(ram_s_70_2), .C(CLK_3P3_MHZ_c), .D(n1450));   // src/ram.vhd(56[12:17])
    SB_DFF i1697_1698 (.Q(ram_s_70_1), .C(CLK_3P3_MHZ_c), .D(n1449));   // src/ram.vhd(56[12:17])
    SB_DFF i1694_1695 (.Q(ram_s_70_0), .C(CLK_3P3_MHZ_c), .D(n1448));   // src/ram.vhd(56[12:17])
    SB_DFF i1691_1692 (.Q(ram_s_69_7), .C(CLK_3P3_MHZ_c), .D(n1447));   // src/ram.vhd(56[12:17])
    SB_DFF i1688_1689 (.Q(ram_s_69_6), .C(CLK_3P3_MHZ_c), .D(n1446));   // src/ram.vhd(56[12:17])
    SB_DFF i1685_1686 (.Q(ram_s_69_5), .C(CLK_3P3_MHZ_c), .D(n1445));   // src/ram.vhd(56[12:17])
    SB_DFF i1682_1683 (.Q(ram_s_69_4), .C(CLK_3P3_MHZ_c), .D(n1444));   // src/ram.vhd(56[12:17])
    SB_DFF i1679_1680 (.Q(ram_s_69_3), .C(CLK_3P3_MHZ_c), .D(n1443));   // src/ram.vhd(56[12:17])
    SB_DFF i1676_1677 (.Q(ram_s_69_2), .C(CLK_3P3_MHZ_c), .D(n1442));   // src/ram.vhd(56[12:17])
    SB_DFF i1673_1674 (.Q(ram_s_69_1), .C(CLK_3P3_MHZ_c), .D(n1441));   // src/ram.vhd(56[12:17])
    SB_DFF i1670_1671 (.Q(ram_s_69_0), .C(CLK_3P3_MHZ_c), .D(n1440));   // src/ram.vhd(56[12:17])
    SB_DFF i1667_1668 (.Q(ram_s_68_7), .C(CLK_3P3_MHZ_c), .D(n1439));   // src/ram.vhd(56[12:17])
    SB_DFF i1664_1665 (.Q(ram_s_68_6), .C(CLK_3P3_MHZ_c), .D(n1438));   // src/ram.vhd(56[12:17])
    SB_DFF i1661_1662 (.Q(ram_s_68_5), .C(CLK_3P3_MHZ_c), .D(n1437));   // src/ram.vhd(56[12:17])
    SB_DFF i1658_1659 (.Q(ram_s_68_4), .C(CLK_3P3_MHZ_c), .D(n1436));   // src/ram.vhd(56[12:17])
    SB_DFF i1655_1656 (.Q(ram_s_68_3), .C(CLK_3P3_MHZ_c), .D(n1435));   // src/ram.vhd(56[12:17])
    SB_DFF i1652_1653 (.Q(ram_s_68_2), .C(CLK_3P3_MHZ_c), .D(n1434));   // src/ram.vhd(56[12:17])
    SB_DFF i1649_1650 (.Q(ram_s_68_1), .C(CLK_3P3_MHZ_c), .D(n1433));   // src/ram.vhd(56[12:17])
    SB_DFF i1646_1647 (.Q(ram_s_68_0), .C(CLK_3P3_MHZ_c), .D(n1432));   // src/ram.vhd(56[12:17])
    SB_DFF i1643_1644 (.Q(ram_s_67_7), .C(CLK_3P3_MHZ_c), .D(n1431));   // src/ram.vhd(56[12:17])
    SB_DFF i1640_1641 (.Q(ram_s_67_6), .C(CLK_3P3_MHZ_c), .D(n1430));   // src/ram.vhd(56[12:17])
    SB_DFF i1637_1638 (.Q(ram_s_67_5), .C(CLK_3P3_MHZ_c), .D(n1429));   // src/ram.vhd(56[12:17])
    SB_DFF i1634_1635 (.Q(ram_s_67_4), .C(CLK_3P3_MHZ_c), .D(n1428));   // src/ram.vhd(56[12:17])
    SB_DFF i1631_1632 (.Q(ram_s_67_3), .C(CLK_3P3_MHZ_c), .D(n1427));   // src/ram.vhd(56[12:17])
    SB_DFF i1628_1629 (.Q(ram_s_67_2), .C(CLK_3P3_MHZ_c), .D(n1426));   // src/ram.vhd(56[12:17])
    SB_DFF i1625_1626 (.Q(ram_s_67_1), .C(CLK_3P3_MHZ_c), .D(n1425));   // src/ram.vhd(56[12:17])
    SB_DFF i1622_1623 (.Q(ram_s_67_0), .C(CLK_3P3_MHZ_c), .D(n1424));   // src/ram.vhd(56[12:17])
    SB_DFF i1619_1620 (.Q(ram_s_66_7), .C(CLK_3P3_MHZ_c), .D(n1423));   // src/ram.vhd(56[12:17])
    SB_DFF i1616_1617 (.Q(ram_s_66_6), .C(CLK_3P3_MHZ_c), .D(n1422));   // src/ram.vhd(56[12:17])
    SB_DFF i1613_1614 (.Q(ram_s_66_5), .C(CLK_3P3_MHZ_c), .D(n1421));   // src/ram.vhd(56[12:17])
    SB_DFF i1610_1611 (.Q(ram_s_66_4), .C(CLK_3P3_MHZ_c), .D(n1420));   // src/ram.vhd(56[12:17])
    SB_DFF i1607_1608 (.Q(ram_s_66_3), .C(CLK_3P3_MHZ_c), .D(n1419));   // src/ram.vhd(56[12:17])
    SB_DFF i1604_1605 (.Q(ram_s_66_2), .C(CLK_3P3_MHZ_c), .D(n1418));   // src/ram.vhd(56[12:17])
    SB_DFF i1601_1602 (.Q(ram_s_66_1), .C(CLK_3P3_MHZ_c), .D(n1417));   // src/ram.vhd(56[12:17])
    SB_DFF i1598_1599 (.Q(ram_s_66_0), .C(CLK_3P3_MHZ_c), .D(n1416));   // src/ram.vhd(56[12:17])
    SB_DFF i1595_1596 (.Q(ram_s_65_7), .C(CLK_3P3_MHZ_c), .D(n1415));   // src/ram.vhd(56[12:17])
    SB_DFF i1592_1593 (.Q(ram_s_65_6), .C(CLK_3P3_MHZ_c), .D(n1414));   // src/ram.vhd(56[12:17])
    SB_DFF i1589_1590 (.Q(ram_s_65_5), .C(CLK_3P3_MHZ_c), .D(n1413));   // src/ram.vhd(56[12:17])
    SB_DFF i1586_1587 (.Q(ram_s_65_4), .C(CLK_3P3_MHZ_c), .D(n1412));   // src/ram.vhd(56[12:17])
    SB_DFF i1583_1584 (.Q(ram_s_65_3), .C(CLK_3P3_MHZ_c), .D(n1411));   // src/ram.vhd(56[12:17])
    SB_DFF i1580_1581 (.Q(ram_s_65_2), .C(CLK_3P3_MHZ_c), .D(n1410));   // src/ram.vhd(56[12:17])
    SB_DFF i1577_1578 (.Q(ram_s_65_1), .C(CLK_3P3_MHZ_c), .D(n1409));   // src/ram.vhd(56[12:17])
    SB_DFF i1574_1575 (.Q(ram_s_65_0), .C(CLK_3P3_MHZ_c), .D(n1408));   // src/ram.vhd(56[12:17])
    SB_DFF i1571_1572 (.Q(ram_s_64_7), .C(CLK_3P3_MHZ_c), .D(n1407));   // src/ram.vhd(56[12:17])
    SB_DFF i1568_1569 (.Q(ram_s_64_6), .C(CLK_3P3_MHZ_c), .D(n1406));   // src/ram.vhd(56[12:17])
    SB_DFF i1565_1566 (.Q(ram_s_64_5), .C(CLK_3P3_MHZ_c), .D(n1405));   // src/ram.vhd(56[12:17])
    SB_DFF i1562_1563 (.Q(ram_s_64_4), .C(CLK_3P3_MHZ_c), .D(n1404));   // src/ram.vhd(56[12:17])
    SB_DFF i1559_1560 (.Q(ram_s_64_3), .C(CLK_3P3_MHZ_c), .D(n1403));   // src/ram.vhd(56[12:17])
    SB_DFF i1556_1557 (.Q(ram_s_64_2), .C(CLK_3P3_MHZ_c), .D(n1402));   // src/ram.vhd(56[12:17])
    SB_DFF i1553_1554 (.Q(ram_s_64_1), .C(CLK_3P3_MHZ_c), .D(n1401));   // src/ram.vhd(56[12:17])
    SB_DFF i1550_1551 (.Q(ram_s_64_0), .C(CLK_3P3_MHZ_c), .D(n1400));   // src/ram.vhd(56[12:17])
    SB_DFF i1547_1548 (.Q(ram_s_63_7), .C(CLK_3P3_MHZ_c), .D(n1399));   // src/ram.vhd(56[12:17])
    SB_DFF i1544_1545 (.Q(ram_s_63_6), .C(CLK_3P3_MHZ_c), .D(n1398));   // src/ram.vhd(56[12:17])
    SB_DFF i1541_1542 (.Q(ram_s_63_5), .C(CLK_3P3_MHZ_c), .D(n1397));   // src/ram.vhd(56[12:17])
    SB_DFF i1538_1539 (.Q(ram_s_63_4), .C(CLK_3P3_MHZ_c), .D(n1396));   // src/ram.vhd(56[12:17])
    SB_DFF i1535_1536 (.Q(ram_s_63_3), .C(CLK_3P3_MHZ_c), .D(n1395));   // src/ram.vhd(56[12:17])
    SB_DFF i1532_1533 (.Q(ram_s_63_2), .C(CLK_3P3_MHZ_c), .D(n1394));   // src/ram.vhd(56[12:17])
    SB_DFF i1529_1530 (.Q(ram_s_63_1), .C(CLK_3P3_MHZ_c), .D(n1393));   // src/ram.vhd(56[12:17])
    SB_DFF i1526_1527 (.Q(ram_s_63_0), .C(CLK_3P3_MHZ_c), .D(n1392));   // src/ram.vhd(56[12:17])
    SB_DFF i1523_1524 (.Q(ram_s_62_7), .C(CLK_3P3_MHZ_c), .D(n1391));   // src/ram.vhd(56[12:17])
    SB_DFF i1520_1521 (.Q(ram_s_62_6), .C(CLK_3P3_MHZ_c), .D(n1390));   // src/ram.vhd(56[12:17])
    SB_DFF i1517_1518 (.Q(ram_s_62_5), .C(CLK_3P3_MHZ_c), .D(n1389));   // src/ram.vhd(56[12:17])
    SB_DFF i1514_1515 (.Q(ram_s_62_4), .C(CLK_3P3_MHZ_c), .D(n1388));   // src/ram.vhd(56[12:17])
    SB_DFF i1511_1512 (.Q(ram_s_62_3), .C(CLK_3P3_MHZ_c), .D(n1387));   // src/ram.vhd(56[12:17])
    SB_DFF i1508_1509 (.Q(ram_s_62_2), .C(CLK_3P3_MHZ_c), .D(n1386));   // src/ram.vhd(56[12:17])
    SB_DFF i1505_1506 (.Q(ram_s_62_1), .C(CLK_3P3_MHZ_c), .D(n1385));   // src/ram.vhd(56[12:17])
    SB_DFF i1502_1503 (.Q(ram_s_62_0), .C(CLK_3P3_MHZ_c), .D(n1384));   // src/ram.vhd(56[12:17])
    SB_DFF i1499_1500 (.Q(ram_s_61_7), .C(CLK_3P3_MHZ_c), .D(n1383));   // src/ram.vhd(56[12:17])
    SB_DFF i1496_1497 (.Q(ram_s_61_6), .C(CLK_3P3_MHZ_c), .D(n1382));   // src/ram.vhd(56[12:17])
    SB_DFF i1493_1494 (.Q(ram_s_61_5), .C(CLK_3P3_MHZ_c), .D(n1381));   // src/ram.vhd(56[12:17])
    SB_DFF i1490_1491 (.Q(ram_s_61_4), .C(CLK_3P3_MHZ_c), .D(n1380));   // src/ram.vhd(56[12:17])
    SB_DFF i1487_1488 (.Q(ram_s_61_3), .C(CLK_3P3_MHZ_c), .D(n1379));   // src/ram.vhd(56[12:17])
    SB_DFF i1484_1485 (.Q(ram_s_61_2), .C(CLK_3P3_MHZ_c), .D(n1378));   // src/ram.vhd(56[12:17])
    SB_DFF i1481_1482 (.Q(ram_s_61_1), .C(CLK_3P3_MHZ_c), .D(n1377));   // src/ram.vhd(56[12:17])
    SB_DFF i1478_1479 (.Q(ram_s_61_0), .C(CLK_3P3_MHZ_c), .D(n1376));   // src/ram.vhd(56[12:17])
    SB_DFF i1475_1476 (.Q(ram_s_60_7), .C(CLK_3P3_MHZ_c), .D(n1375));   // src/ram.vhd(56[12:17])
    SB_DFF i1472_1473 (.Q(ram_s_60_6), .C(CLK_3P3_MHZ_c), .D(n1374));   // src/ram.vhd(56[12:17])
    SB_DFF i1469_1470 (.Q(ram_s_60_5), .C(CLK_3P3_MHZ_c), .D(n1373));   // src/ram.vhd(56[12:17])
    SB_DFF i1466_1467 (.Q(ram_s_60_4), .C(CLK_3P3_MHZ_c), .D(n1372));   // src/ram.vhd(56[12:17])
    SB_DFF i1463_1464 (.Q(ram_s_60_3), .C(CLK_3P3_MHZ_c), .D(n1371));   // src/ram.vhd(56[12:17])
    SB_DFF i1460_1461 (.Q(ram_s_60_2), .C(CLK_3P3_MHZ_c), .D(n1370));   // src/ram.vhd(56[12:17])
    SB_DFF i1457_1458 (.Q(ram_s_60_1), .C(CLK_3P3_MHZ_c), .D(n1369));   // src/ram.vhd(56[12:17])
    SB_DFF i1454_1455 (.Q(ram_s_60_0), .C(CLK_3P3_MHZ_c), .D(n1368));   // src/ram.vhd(56[12:17])
    SB_DFF i1451_1452 (.Q(ram_s_59_7), .C(CLK_3P3_MHZ_c), .D(n1367));   // src/ram.vhd(56[12:17])
    SB_DFF i1448_1449 (.Q(ram_s_59_6), .C(CLK_3P3_MHZ_c), .D(n1366));   // src/ram.vhd(56[12:17])
    SB_DFF i1445_1446 (.Q(ram_s_59_5), .C(CLK_3P3_MHZ_c), .D(n1365));   // src/ram.vhd(56[12:17])
    SB_DFF i1442_1443 (.Q(ram_s_59_4), .C(CLK_3P3_MHZ_c), .D(n1364));   // src/ram.vhd(56[12:17])
    SB_DFF i1439_1440 (.Q(ram_s_59_3), .C(CLK_3P3_MHZ_c), .D(n1363));   // src/ram.vhd(56[12:17])
    SB_DFF i1436_1437 (.Q(ram_s_59_2), .C(CLK_3P3_MHZ_c), .D(n1362));   // src/ram.vhd(56[12:17])
    SB_DFF i1433_1434 (.Q(ram_s_59_1), .C(CLK_3P3_MHZ_c), .D(n1361));   // src/ram.vhd(56[12:17])
    SB_DFF i1430_1431 (.Q(ram_s_59_0), .C(CLK_3P3_MHZ_c), .D(n1360));   // src/ram.vhd(56[12:17])
    SB_DFF i1427_1428 (.Q(ram_s_58_7), .C(CLK_3P3_MHZ_c), .D(n1359));   // src/ram.vhd(56[12:17])
    SB_DFF i1424_1425 (.Q(ram_s_58_6), .C(CLK_3P3_MHZ_c), .D(n1358));   // src/ram.vhd(56[12:17])
    SB_DFF i1421_1422 (.Q(ram_s_58_5), .C(CLK_3P3_MHZ_c), .D(n1357));   // src/ram.vhd(56[12:17])
    SB_DFF i1418_1419 (.Q(ram_s_58_4), .C(CLK_3P3_MHZ_c), .D(n1356));   // src/ram.vhd(56[12:17])
    SB_DFF i1415_1416 (.Q(ram_s_58_3), .C(CLK_3P3_MHZ_c), .D(n1355));   // src/ram.vhd(56[12:17])
    SB_DFF i1412_1413 (.Q(ram_s_58_2), .C(CLK_3P3_MHZ_c), .D(n1354));   // src/ram.vhd(56[12:17])
    SB_DFF i1409_1410 (.Q(ram_s_58_1), .C(CLK_3P3_MHZ_c), .D(n1353));   // src/ram.vhd(56[12:17])
    SB_DFF i1406_1407 (.Q(ram_s_58_0), .C(CLK_3P3_MHZ_c), .D(n1352));   // src/ram.vhd(56[12:17])
    SB_DFF i1403_1404 (.Q(ram_s_57_7), .C(CLK_3P3_MHZ_c), .D(n1351));   // src/ram.vhd(56[12:17])
    SB_DFF i1400_1401 (.Q(ram_s_57_6), .C(CLK_3P3_MHZ_c), .D(n1350));   // src/ram.vhd(56[12:17])
    SB_DFF i1397_1398 (.Q(ram_s_57_5), .C(CLK_3P3_MHZ_c), .D(n1349));   // src/ram.vhd(56[12:17])
    SB_DFF i1394_1395 (.Q(ram_s_57_4), .C(CLK_3P3_MHZ_c), .D(n1348));   // src/ram.vhd(56[12:17])
    SB_DFF i1391_1392 (.Q(ram_s_57_3), .C(CLK_3P3_MHZ_c), .D(n1347));   // src/ram.vhd(56[12:17])
    SB_DFF i1388_1389 (.Q(ram_s_57_2), .C(CLK_3P3_MHZ_c), .D(n1346));   // src/ram.vhd(56[12:17])
    SB_DFF i1385_1386 (.Q(ram_s_57_1), .C(CLK_3P3_MHZ_c), .D(n1345));   // src/ram.vhd(56[12:17])
    SB_DFF i1382_1383 (.Q(ram_s_57_0), .C(CLK_3P3_MHZ_c), .D(n1344));   // src/ram.vhd(56[12:17])
    SB_DFF i1379_1380 (.Q(ram_s_56_7), .C(CLK_3P3_MHZ_c), .D(n1343));   // src/ram.vhd(56[12:17])
    SB_DFF i1376_1377 (.Q(ram_s_56_6), .C(CLK_3P3_MHZ_c), .D(n1342));   // src/ram.vhd(56[12:17])
    SB_DFF i1373_1374 (.Q(ram_s_56_5), .C(CLK_3P3_MHZ_c), .D(n1341));   // src/ram.vhd(56[12:17])
    SB_DFF i1370_1371 (.Q(ram_s_56_4), .C(CLK_3P3_MHZ_c), .D(n1340));   // src/ram.vhd(56[12:17])
    SB_DFF i1367_1368 (.Q(ram_s_56_3), .C(CLK_3P3_MHZ_c), .D(n1339));   // src/ram.vhd(56[12:17])
    SB_DFF i1364_1365 (.Q(ram_s_56_2), .C(CLK_3P3_MHZ_c), .D(n1338));   // src/ram.vhd(56[12:17])
    SB_DFF i1361_1362 (.Q(ram_s_56_1), .C(CLK_3P3_MHZ_c), .D(n1337));   // src/ram.vhd(56[12:17])
    SB_DFF i1358_1359 (.Q(ram_s_56_0), .C(CLK_3P3_MHZ_c), .D(n1336));   // src/ram.vhd(56[12:17])
    SB_DFF i1355_1356 (.Q(ram_s_55_7), .C(CLK_3P3_MHZ_c), .D(n1335));   // src/ram.vhd(56[12:17])
    SB_DFF i1352_1353 (.Q(ram_s_55_6), .C(CLK_3P3_MHZ_c), .D(n1334));   // src/ram.vhd(56[12:17])
    SB_DFF i1349_1350 (.Q(ram_s_55_5), .C(CLK_3P3_MHZ_c), .D(n1333));   // src/ram.vhd(56[12:17])
    SB_DFF i1346_1347 (.Q(ram_s_55_4), .C(CLK_3P3_MHZ_c), .D(n1332));   // src/ram.vhd(56[12:17])
    SB_DFF i1343_1344 (.Q(ram_s_55_3), .C(CLK_3P3_MHZ_c), .D(n1331));   // src/ram.vhd(56[12:17])
    SB_DFF i1340_1341 (.Q(ram_s_55_2), .C(CLK_3P3_MHZ_c), .D(n1330));   // src/ram.vhd(56[12:17])
    SB_DFF i1337_1338 (.Q(ram_s_55_1), .C(CLK_3P3_MHZ_c), .D(n1329));   // src/ram.vhd(56[12:17])
    SB_DFF i1334_1335 (.Q(ram_s_55_0), .C(CLK_3P3_MHZ_c), .D(n1328));   // src/ram.vhd(56[12:17])
    SB_DFF i1331_1332 (.Q(ram_s_54_7), .C(CLK_3P3_MHZ_c), .D(n1327));   // src/ram.vhd(56[12:17])
    SB_DFF i1328_1329 (.Q(ram_s_54_6), .C(CLK_3P3_MHZ_c), .D(n1326));   // src/ram.vhd(56[12:17])
    SB_DFF i1325_1326 (.Q(ram_s_54_5), .C(CLK_3P3_MHZ_c), .D(n1325));   // src/ram.vhd(56[12:17])
    SB_DFF i1322_1323 (.Q(ram_s_54_4), .C(CLK_3P3_MHZ_c), .D(n1324));   // src/ram.vhd(56[12:17])
    SB_DFF i1319_1320 (.Q(ram_s_54_3), .C(CLK_3P3_MHZ_c), .D(n1323));   // src/ram.vhd(56[12:17])
    SB_DFF i1316_1317 (.Q(ram_s_54_2), .C(CLK_3P3_MHZ_c), .D(n1322));   // src/ram.vhd(56[12:17])
    SB_DFF i1313_1314 (.Q(ram_s_54_1), .C(CLK_3P3_MHZ_c), .D(n1321));   // src/ram.vhd(56[12:17])
    SB_DFF i1310_1311 (.Q(ram_s_54_0), .C(CLK_3P3_MHZ_c), .D(n1320));   // src/ram.vhd(56[12:17])
    SB_DFF i1307_1308 (.Q(ram_s_53_7), .C(CLK_3P3_MHZ_c), .D(n1319));   // src/ram.vhd(56[12:17])
    SB_DFF i1304_1305 (.Q(ram_s_53_6), .C(CLK_3P3_MHZ_c), .D(n1318));   // src/ram.vhd(56[12:17])
    SB_DFF i1301_1302 (.Q(ram_s_53_5), .C(CLK_3P3_MHZ_c), .D(n1317));   // src/ram.vhd(56[12:17])
    SB_DFF i1298_1299 (.Q(ram_s_53_4), .C(CLK_3P3_MHZ_c), .D(n1316));   // src/ram.vhd(56[12:17])
    SB_DFF i1295_1296 (.Q(ram_s_53_3), .C(CLK_3P3_MHZ_c), .D(n1315));   // src/ram.vhd(56[12:17])
    SB_DFF i1292_1293 (.Q(ram_s_53_2), .C(CLK_3P3_MHZ_c), .D(n1314));   // src/ram.vhd(56[12:17])
    SB_DFF i1289_1290 (.Q(ram_s_53_1), .C(CLK_3P3_MHZ_c), .D(n1313));   // src/ram.vhd(56[12:17])
    SB_DFF i1286_1287 (.Q(ram_s_53_0), .C(CLK_3P3_MHZ_c), .D(n1312));   // src/ram.vhd(56[12:17])
    SB_DFF i1283_1284 (.Q(ram_s_52_7), .C(CLK_3P3_MHZ_c), .D(n1311));   // src/ram.vhd(56[12:17])
    SB_DFF i1280_1281 (.Q(ram_s_52_6), .C(CLK_3P3_MHZ_c), .D(n1310));   // src/ram.vhd(56[12:17])
    SB_DFF i1277_1278 (.Q(ram_s_52_5), .C(CLK_3P3_MHZ_c), .D(n1309));   // src/ram.vhd(56[12:17])
    SB_DFF i1274_1275 (.Q(ram_s_52_4), .C(CLK_3P3_MHZ_c), .D(n1308));   // src/ram.vhd(56[12:17])
    SB_DFF i1271_1272 (.Q(ram_s_52_3), .C(CLK_3P3_MHZ_c), .D(n1307));   // src/ram.vhd(56[12:17])
    SB_DFF i1268_1269 (.Q(ram_s_52_2), .C(CLK_3P3_MHZ_c), .D(n1306));   // src/ram.vhd(56[12:17])
    SB_DFF i1265_1266 (.Q(ram_s_52_1), .C(CLK_3P3_MHZ_c), .D(n1305));   // src/ram.vhd(56[12:17])
    SB_DFF i1262_1263 (.Q(ram_s_52_0), .C(CLK_3P3_MHZ_c), .D(n1304));   // src/ram.vhd(56[12:17])
    SB_DFF i1259_1260 (.Q(ram_s_51_7), .C(CLK_3P3_MHZ_c), .D(n1303));   // src/ram.vhd(56[12:17])
    SB_DFF i1256_1257 (.Q(ram_s_51_6), .C(CLK_3P3_MHZ_c), .D(n1302));   // src/ram.vhd(56[12:17])
    SB_DFF i1253_1254 (.Q(ram_s_51_5), .C(CLK_3P3_MHZ_c), .D(n1301));   // src/ram.vhd(56[12:17])
    SB_LUT4 i707_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_20_0), .O(n955));   // src/ram.vhd(68[19:45])
    defparam i707_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1250_1251 (.Q(ram_s_51_4), .C(CLK_3P3_MHZ_c), .D(n1300));   // src/ram.vhd(56[12:17])
    SB_LUT4 i674_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_20_7), .O(n922));   // src/ram.vhd(68[19:45])
    defparam i674_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1247_1248 (.Q(ram_s_51_3), .C(CLK_3P3_MHZ_c), .D(n1299));   // src/ram.vhd(56[12:17])
    SB_LUT4 i681_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_20_6), .O(n929));   // src/ram.vhd(68[19:45])
    defparam i681_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1244_1245 (.Q(ram_s_51_2), .C(CLK_3P3_MHZ_c), .D(n1298));   // src/ram.vhd(56[12:17])
    SB_LUT4 i694_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_20_5), .O(n942));   // src/ram.vhd(68[19:45])
    defparam i694_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1241_1242 (.Q(ram_s_51_1), .C(CLK_3P3_MHZ_c), .D(n1297));   // src/ram.vhd(56[12:17])
    SB_LUT4 i695_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_20_4), .O(n943));   // src/ram.vhd(68[19:45])
    defparam i695_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1238_1239 (.Q(ram_s_51_0), .C(CLK_3P3_MHZ_c), .D(n1296));   // src/ram.vhd(56[12:17])
    SB_LUT4 i697_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_20_3), .O(n945));   // src/ram.vhd(68[19:45])
    defparam i697_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1235_1236 (.Q(ram_s_50_7), .C(CLK_3P3_MHZ_c), .D(n1295));   // src/ram.vhd(56[12:17])
    SB_LUT4 i699_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_20_2), .O(n947));   // src/ram.vhd(68[19:45])
    defparam i699_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1232_1233 (.Q(ram_s_50_6), .C(CLK_3P3_MHZ_c), .D(n1294));   // src/ram.vhd(56[12:17])
    SB_LUT4 i706_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_20_1), .O(n954));   // src/ram.vhd(68[19:45])
    defparam i706_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1229_1230 (.Q(ram_s_50_5), .C(CLK_3P3_MHZ_c), .D(n1293));   // src/ram.vhd(56[12:17])
    SB_LUT4 i776_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_18_2), .O(n1024));   // src/ram.vhd(68[19:45])
    defparam i776_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1226_1227 (.Q(ram_s_50_4), .C(CLK_3P3_MHZ_c), .D(n1292));   // src/ram.vhd(56[12:17])
    SB_LUT4 i772_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_18_6), .O(n1020));   // src/ram.vhd(68[19:45])
    defparam i772_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1223_1224 (.Q(ram_s_50_3), .C(CLK_3P3_MHZ_c), .D(n1291));   // src/ram.vhd(56[12:17])
    SB_LUT4 i773_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_18_5), .O(n1021));   // src/ram.vhd(68[19:45])
    defparam i773_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1220_1221 (.Q(ram_s_50_2), .C(CLK_3P3_MHZ_c), .D(n1290));   // src/ram.vhd(56[12:17])
    SB_LUT4 i774_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_18_4), .O(n1022));   // src/ram.vhd(68[19:45])
    defparam i774_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1217_1218 (.Q(ram_s_50_1), .C(CLK_3P3_MHZ_c), .D(n1289));   // src/ram.vhd(56[12:17])
    SB_LUT4 i775_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_18_3), .O(n1023));   // src/ram.vhd(68[19:45])
    defparam i775_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1214_1215 (.Q(ram_s_50_0), .C(CLK_3P3_MHZ_c), .D(n1288));   // src/ram.vhd(56[12:17])
    SB_LUT4 i771_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_18_7), .O(n1019));   // src/ram.vhd(68[19:45])
    defparam i771_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1211_1212 (.Q(ram_s_49_7), .C(CLK_3P3_MHZ_c), .D(n1287));   // src/ram.vhd(56[12:17])
    SB_LUT4 i671_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_18_1), .O(n919));   // src/ram.vhd(68[19:45])
    defparam i671_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1208_1209 (.Q(ram_s_49_6), .C(CLK_3P3_MHZ_c), .D(n1286));   // src/ram.vhd(56[12:17])
    SB_LUT4 i673_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_18_0), .O(n921));   // src/ram.vhd(68[19:45])
    defparam i673_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1205_1206 (.Q(ram_s_49_5), .C(CLK_3P3_MHZ_c), .D(n1285));   // src/ram.vhd(56[12:17])
    SB_LUT4 i809_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_19_2), .O(n1057));   // src/ram.vhd(68[19:45])
    defparam i809_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1202_1203 (.Q(ram_s_49_4), .C(CLK_3P3_MHZ_c), .D(n1284));   // src/ram.vhd(56[12:17])
    SB_LUT4 i779_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_19_5), .O(n1027));   // src/ram.vhd(68[19:45])
    defparam i779_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1199_1200 (.Q(ram_s_49_3), .C(CLK_3P3_MHZ_c), .D(n1283));   // src/ram.vhd(56[12:17])
    SB_LUT4 i780_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_19_4), .O(n1028));   // src/ram.vhd(68[19:45])
    defparam i780_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1196_1197 (.Q(ram_s_49_2), .C(CLK_3P3_MHZ_c), .D(n1282));   // src/ram.vhd(56[12:17])
    SB_LUT4 i802_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_19_3), .O(n1050));   // src/ram.vhd(68[19:45])
    defparam i802_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1193_1194 (.Q(ram_s_49_1), .C(CLK_3P3_MHZ_c), .D(n1281));   // src/ram.vhd(56[12:17])
    SB_LUT4 i666_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_19_1), .O(n914));   // src/ram.vhd(68[19:45])
    defparam i666_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1190_1191 (.Q(ram_s_49_0), .C(CLK_3P3_MHZ_c), .D(n1280));   // src/ram.vhd(56[12:17])
    SB_LUT4 i770_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_19_0), .O(n1018));   // src/ram.vhd(68[19:45])
    defparam i770_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1187_1188 (.Q(ram_s_48_7), .C(CLK_3P3_MHZ_c), .D(n1279));   // src/ram.vhd(56[12:17])
    SB_LUT4 i777_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_19_7), .O(n1025));   // src/ram.vhd(68[19:45])
    defparam i777_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1184_1185 (.Q(ram_s_48_6), .C(CLK_3P3_MHZ_c), .D(n1278));   // src/ram.vhd(56[12:17])
    SB_LUT4 i778_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_19_6), .O(n1026));   // src/ram.vhd(68[19:45])
    defparam i778_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1181_1182 (.Q(ram_s_48_5), .C(CLK_3P3_MHZ_c), .D(n1277));   // src/ram.vhd(56[12:17])
    SB_LUT4 i811_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_16_0), .O(n1059));   // src/ram.vhd(68[19:45])
    defparam i811_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1178_1179 (.Q(ram_s_48_4), .C(CLK_3P3_MHZ_c), .D(n1276));   // src/ram.vhd(56[12:17])
    SB_LUT4 i703_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_16_7), .O(n951));   // src/ram.vhd(68[19:45])
    defparam i703_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1175_1176 (.Q(ram_s_48_3), .C(CLK_3P3_MHZ_c), .D(n1275));   // src/ram.vhd(56[12:17])
    SB_LUT4 i705_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_16_6), .O(n953));   // src/ram.vhd(68[19:45])
    defparam i705_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1172_1173 (.Q(ram_s_48_2), .C(CLK_3P3_MHZ_c), .D(n1274));   // src/ram.vhd(56[12:17])
    SB_LUT4 i800_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_16_5), .O(n1048));   // src/ram.vhd(68[19:45])
    defparam i800_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1169_1170 (.Q(ram_s_48_1), .C(CLK_3P3_MHZ_c), .D(n1273));   // src/ram.vhd(56[12:17])
    SB_LUT4 i805_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_16_4), .O(n1053));   // src/ram.vhd(68[19:45])
    defparam i805_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1166_1167 (.Q(ram_s_48_0), .C(CLK_3P3_MHZ_c), .D(n1272));   // src/ram.vhd(56[12:17])
    SB_LUT4 i806_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_16_3), .O(n1054));   // src/ram.vhd(68[19:45])
    defparam i806_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1163_1164 (.Q(ram_s_47_7), .C(CLK_3P3_MHZ_c), .D(n1271));   // src/ram.vhd(56[12:17])
    SB_LUT4 i807_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_16_2), .O(n1055));   // src/ram.vhd(68[19:45])
    defparam i807_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1160_1161 (.Q(ram_s_47_6), .C(CLK_3P3_MHZ_c), .D(n1270));   // src/ram.vhd(56[12:17])
    SB_LUT4 i810_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_16_1), .O(n1058));   // src/ram.vhd(68[19:45])
    defparam i810_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1157_1158 (.Q(ram_s_47_5), .C(CLK_3P3_MHZ_c), .D(n1269));   // src/ram.vhd(56[12:17])
    SB_LUT4 i812_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_15_7), .O(n1060));   // src/ram.vhd(68[19:45])
    defparam i812_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1154_1155 (.Q(ram_s_47_4), .C(CLK_3P3_MHZ_c), .D(n1268));   // src/ram.vhd(56[12:17])
    SB_LUT4 i652_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_15_4), .O(n900));   // src/ram.vhd(68[19:45])
    defparam i652_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1151_1152 (.Q(ram_s_47_3), .C(CLK_3P3_MHZ_c), .D(n1267));   // src/ram.vhd(56[12:17])
    SB_LUT4 i654_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_15_3), .O(n902));   // src/ram.vhd(68[19:45])
    defparam i654_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1148_1149 (.Q(ram_s_47_2), .C(CLK_3P3_MHZ_c), .D(n1266));   // src/ram.vhd(56[12:17])
    SB_LUT4 i655_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_15_2), .O(n903));   // src/ram.vhd(68[19:45])
    defparam i655_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1145_1146 (.Q(ram_s_47_1), .C(CLK_3P3_MHZ_c), .D(n1265));   // src/ram.vhd(56[12:17])
    SB_LUT4 i665_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_15_1), .O(n913));   // src/ram.vhd(68[19:45])
    defparam i665_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1142_1143 (.Q(ram_s_47_0), .C(CLK_3P3_MHZ_c), .D(n1264));   // src/ram.vhd(56[12:17])
    SB_LUT4 i708_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_15_0), .O(n956));   // src/ram.vhd(68[19:45])
    defparam i708_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1139_1140 (.Q(ram_s_46_7), .C(CLK_3P3_MHZ_c), .D(n1263));   // src/ram.vhd(56[12:17])
    SB_LUT4 i801_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_15_6), .O(n1049));   // src/ram.vhd(68[19:45])
    defparam i801_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1136_1137 (.Q(ram_s_46_6), .C(CLK_3P3_MHZ_c), .D(n1262));   // src/ram.vhd(56[12:17])
    SB_LUT4 i804_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_15_5), .O(n1052));   // src/ram.vhd(68[19:45])
    defparam i804_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1133_1134 (.Q(ram_s_46_5), .C(CLK_3P3_MHZ_c), .D(n1261));   // src/ram.vhd(56[12:17])
    SB_LUT4 i823_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_22_7), .O(n1071));   // src/ram.vhd(68[19:45])
    defparam i823_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1130_1131 (.Q(ram_s_46_4), .C(CLK_3P3_MHZ_c), .D(n1260));   // src/ram.vhd(56[12:17])
    SB_LUT4 i822_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_22_6), .O(n1070));   // src/ram.vhd(68[19:45])
    defparam i822_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1127_1128 (.Q(ram_s_46_3), .C(CLK_3P3_MHZ_c), .D(n1259));   // src/ram.vhd(56[12:17])
    SB_LUT4 i821_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_22_5), .O(n1069));   // src/ram.vhd(68[19:45])
    defparam i821_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1124_1125 (.Q(ram_s_46_2), .C(CLK_3P3_MHZ_c), .D(n1258));   // src/ram.vhd(56[12:17])
    SB_LUT4 i820_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_22_4), .O(n1068));   // src/ram.vhd(68[19:45])
    defparam i820_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1121_1122 (.Q(ram_s_46_1), .C(CLK_3P3_MHZ_c), .D(n1257));   // src/ram.vhd(56[12:17])
    SB_LUT4 i819_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_22_3), .O(n1067));   // src/ram.vhd(68[19:45])
    defparam i819_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1118_1119 (.Q(ram_s_46_0), .C(CLK_3P3_MHZ_c), .D(n1256));   // src/ram.vhd(56[12:17])
    SB_LUT4 i818_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_22_2), .O(n1066));   // src/ram.vhd(68[19:45])
    defparam i818_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1115_1116 (.Q(ram_s_45_7), .C(CLK_3P3_MHZ_c), .D(n1255));   // src/ram.vhd(56[12:17])
    SB_LUT4 i817_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_22_1), .O(n1065));   // src/ram.vhd(68[19:45])
    defparam i817_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1112_1113 (.Q(ram_s_45_6), .C(CLK_3P3_MHZ_c), .D(n1254));   // src/ram.vhd(56[12:17])
    SB_LUT4 i816_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_22_0), .O(n1064));   // src/ram.vhd(68[19:45])
    defparam i816_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1109_1110 (.Q(ram_s_45_5), .C(CLK_3P3_MHZ_c), .D(n1253));   // src/ram.vhd(56[12:17])
    SB_LUT4 i831_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_23_7), .O(n1079));   // src/ram.vhd(68[19:45])
    defparam i831_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1106_1107 (.Q(ram_s_45_4), .C(CLK_3P3_MHZ_c), .D(n1252));   // src/ram.vhd(56[12:17])
    SB_LUT4 i830_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_23_6), .O(n1078));   // src/ram.vhd(68[19:45])
    defparam i830_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1103_1104 (.Q(ram_s_45_3), .C(CLK_3P3_MHZ_c), .D(n1251));   // src/ram.vhd(56[12:17])
    SB_LUT4 i829_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_23_5), .O(n1077));   // src/ram.vhd(68[19:45])
    defparam i829_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1100_1101 (.Q(ram_s_45_2), .C(CLK_3P3_MHZ_c), .D(n1250));   // src/ram.vhd(56[12:17])
    SB_LUT4 i828_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_23_4), .O(n1076));   // src/ram.vhd(68[19:45])
    defparam i828_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1097_1098 (.Q(ram_s_45_1), .C(CLK_3P3_MHZ_c), .D(n1249));   // src/ram.vhd(56[12:17])
    SB_LUT4 i827_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_23_3), .O(n1075));   // src/ram.vhd(68[19:45])
    defparam i827_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1094_1095 (.Q(ram_s_45_0), .C(CLK_3P3_MHZ_c), .D(n1248));   // src/ram.vhd(56[12:17])
    SB_LUT4 i826_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_23_2), .O(n1074));   // src/ram.vhd(68[19:45])
    defparam i826_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1091_1092 (.Q(ram_s_44_7), .C(CLK_3P3_MHZ_c), .D(n1247));   // src/ram.vhd(56[12:17])
    SB_LUT4 i825_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_23_1), .O(n1073));   // src/ram.vhd(68[19:45])
    defparam i825_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1088_1089 (.Q(ram_s_44_6), .C(CLK_3P3_MHZ_c), .D(n1246));   // src/ram.vhd(56[12:17])
    SB_LUT4 i824_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_23_0), .O(n1072));   // src/ram.vhd(68[19:45])
    defparam i824_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1085_1086 (.Q(ram_s_44_5), .C(CLK_3P3_MHZ_c), .D(n1245));   // src/ram.vhd(56[12:17])
    SB_LUT4 i839_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_24_7), .O(n1087));   // src/ram.vhd(68[19:45])
    defparam i839_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1082_1083 (.Q(ram_s_44_4), .C(CLK_3P3_MHZ_c), .D(n1244));   // src/ram.vhd(56[12:17])
    SB_LUT4 i838_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_24_6), .O(n1086));   // src/ram.vhd(68[19:45])
    defparam i838_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1079_1080 (.Q(ram_s_44_3), .C(CLK_3P3_MHZ_c), .D(n1243));   // src/ram.vhd(56[12:17])
    SB_LUT4 i837_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_24_5), .O(n1085));   // src/ram.vhd(68[19:45])
    defparam i837_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1076_1077 (.Q(ram_s_44_2), .C(CLK_3P3_MHZ_c), .D(n1242));   // src/ram.vhd(56[12:17])
    SB_LUT4 i836_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_24_4), .O(n1084));   // src/ram.vhd(68[19:45])
    defparam i836_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1073_1074 (.Q(ram_s_44_1), .C(CLK_3P3_MHZ_c), .D(n1241));   // src/ram.vhd(56[12:17])
    SB_LUT4 i835_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_24_3), .O(n1083));   // src/ram.vhd(68[19:45])
    defparam i835_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1070_1071 (.Q(ram_s_44_0), .C(CLK_3P3_MHZ_c), .D(n1240));   // src/ram.vhd(56[12:17])
    SB_LUT4 i834_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_24_2), .O(n1082));   // src/ram.vhd(68[19:45])
    defparam i834_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1067_1068 (.Q(ram_s_43_7), .C(CLK_3P3_MHZ_c), .D(n1239));   // src/ram.vhd(56[12:17])
    SB_LUT4 i833_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_24_1), .O(n1081));   // src/ram.vhd(68[19:45])
    defparam i833_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1064_1065 (.Q(ram_s_43_6), .C(CLK_3P3_MHZ_c), .D(n1238));   // src/ram.vhd(56[12:17])
    SB_LUT4 i832_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_24_0), .O(n1080));   // src/ram.vhd(68[19:45])
    defparam i832_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1061_1062 (.Q(ram_s_43_5), .C(CLK_3P3_MHZ_c), .D(n1237));   // src/ram.vhd(56[12:17])
    SB_LUT4 i847_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_25_7), .O(n1095));   // src/ram.vhd(68[19:45])
    defparam i847_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1058_1059 (.Q(ram_s_43_4), .C(CLK_3P3_MHZ_c), .D(n1236));   // src/ram.vhd(56[12:17])
    SB_LUT4 i846_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_25_6), .O(n1094));   // src/ram.vhd(68[19:45])
    defparam i846_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1055_1056 (.Q(ram_s_43_3), .C(CLK_3P3_MHZ_c), .D(n1235));   // src/ram.vhd(56[12:17])
    SB_LUT4 i845_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_25_5), .O(n1093));   // src/ram.vhd(68[19:45])
    defparam i845_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1052_1053 (.Q(ram_s_43_2), .C(CLK_3P3_MHZ_c), .D(n1234));   // src/ram.vhd(56[12:17])
    SB_LUT4 i844_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_25_4), .O(n1092));   // src/ram.vhd(68[19:45])
    defparam i844_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1049_1050 (.Q(ram_s_43_1), .C(CLK_3P3_MHZ_c), .D(n1233));   // src/ram.vhd(56[12:17])
    SB_LUT4 i843_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_25_3), .O(n1091));   // src/ram.vhd(68[19:45])
    defparam i843_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1046_1047 (.Q(ram_s_43_0), .C(CLK_3P3_MHZ_c), .D(n1232));   // src/ram.vhd(56[12:17])
    SB_LUT4 i842_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_25_2), .O(n1090));   // src/ram.vhd(68[19:45])
    defparam i842_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1043_1044 (.Q(ram_s_42_7), .C(CLK_3P3_MHZ_c), .D(n1231));   // src/ram.vhd(56[12:17])
    SB_LUT4 i841_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_25_1), .O(n1089));   // src/ram.vhd(68[19:45])
    defparam i841_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1040_1041 (.Q(ram_s_42_6), .C(CLK_3P3_MHZ_c), .D(n1230));   // src/ram.vhd(56[12:17])
    SB_LUT4 i840_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_25_0), .O(n1088));   // src/ram.vhd(68[19:45])
    defparam i840_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1037_1038 (.Q(ram_s_42_5), .C(CLK_3P3_MHZ_c), .D(n1229));   // src/ram.vhd(56[12:17])
    SB_LUT4 i855_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_26_7), .O(n1103));   // src/ram.vhd(68[19:45])
    defparam i855_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1034_1035 (.Q(ram_s_42_4), .C(CLK_3P3_MHZ_c), .D(n1228));   // src/ram.vhd(56[12:17])
    SB_LUT4 i854_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_26_6), .O(n1102));   // src/ram.vhd(68[19:45])
    defparam i854_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1031_1032 (.Q(ram_s_42_3), .C(CLK_3P3_MHZ_c), .D(n1227));   // src/ram.vhd(56[12:17])
    SB_LUT4 i853_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_26_5), .O(n1101));   // src/ram.vhd(68[19:45])
    defparam i853_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1028_1029 (.Q(ram_s_42_2), .C(CLK_3P3_MHZ_c), .D(n1226));   // src/ram.vhd(56[12:17])
    SB_LUT4 i852_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_26_4), .O(n1100));   // src/ram.vhd(68[19:45])
    defparam i852_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1025_1026 (.Q(ram_s_42_1), .C(CLK_3P3_MHZ_c), .D(n1225));   // src/ram.vhd(56[12:17])
    SB_LUT4 i851_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_26_3), .O(n1099));   // src/ram.vhd(68[19:45])
    defparam i851_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1022_1023 (.Q(ram_s_42_0), .C(CLK_3P3_MHZ_c), .D(n1224));   // src/ram.vhd(56[12:17])
    SB_LUT4 i850_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_26_2), .O(n1098));   // src/ram.vhd(68[19:45])
    defparam i850_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1019_1020 (.Q(ram_s_41_7), .C(CLK_3P3_MHZ_c), .D(n1223));   // src/ram.vhd(56[12:17])
    SB_LUT4 i849_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_26_1), .O(n1097));   // src/ram.vhd(68[19:45])
    defparam i849_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1016_1017 (.Q(ram_s_41_6), .C(CLK_3P3_MHZ_c), .D(n1222));   // src/ram.vhd(56[12:17])
    SB_LUT4 i848_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_26_0), .O(n1096));   // src/ram.vhd(68[19:45])
    defparam i848_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1013_1014 (.Q(ram_s_41_5), .C(CLK_3P3_MHZ_c), .D(n1221));   // src/ram.vhd(56[12:17])
    SB_LUT4 i863_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_27_7), .O(n1111));   // src/ram.vhd(68[19:45])
    defparam i863_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1010_1011 (.Q(ram_s_41_4), .C(CLK_3P3_MHZ_c), .D(n1220));   // src/ram.vhd(56[12:17])
    SB_LUT4 i862_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_27_6), .O(n1110));   // src/ram.vhd(68[19:45])
    defparam i862_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1007_1008 (.Q(ram_s_41_3), .C(CLK_3P3_MHZ_c), .D(n1219));   // src/ram.vhd(56[12:17])
    SB_LUT4 i861_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_27_5), .O(n1109));   // src/ram.vhd(68[19:45])
    defparam i861_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1004_1005 (.Q(ram_s_41_2), .C(CLK_3P3_MHZ_c), .D(n1218));   // src/ram.vhd(56[12:17])
    SB_LUT4 i860_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_27_4), .O(n1108));   // src/ram.vhd(68[19:45])
    defparam i860_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1001_1002 (.Q(ram_s_41_1), .C(CLK_3P3_MHZ_c), .D(n1217));   // src/ram.vhd(56[12:17])
    SB_LUT4 i859_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_27_3), .O(n1107));   // src/ram.vhd(68[19:45])
    defparam i859_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i998_999 (.Q(ram_s_41_0), .C(CLK_3P3_MHZ_c), .D(n1216));   // src/ram.vhd(56[12:17])
    SB_LUT4 i858_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_27_2), .O(n1106));   // src/ram.vhd(68[19:45])
    defparam i858_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i995_996 (.Q(ram_s_40_7), .C(CLK_3P3_MHZ_c), .D(n1215));   // src/ram.vhd(56[12:17])
    SB_LUT4 i857_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_27_1), .O(n1105));   // src/ram.vhd(68[19:45])
    defparam i857_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i992_993 (.Q(ram_s_40_6), .C(CLK_3P3_MHZ_c), .D(n1214));   // src/ram.vhd(56[12:17])
    SB_LUT4 i856_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_27_0), .O(n1104));   // src/ram.vhd(68[19:45])
    defparam i856_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i989_990 (.Q(ram_s_40_5), .C(CLK_3P3_MHZ_c), .D(n1213));   // src/ram.vhd(56[12:17])
    SB_LUT4 i871_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_28_7), .O(n1119));   // src/ram.vhd(68[19:45])
    defparam i871_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i986_987 (.Q(ram_s_40_4), .C(CLK_3P3_MHZ_c), .D(n1212));   // src/ram.vhd(56[12:17])
    SB_LUT4 i870_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_28_6), .O(n1118));   // src/ram.vhd(68[19:45])
    defparam i870_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i983_984 (.Q(ram_s_40_3), .C(CLK_3P3_MHZ_c), .D(n1211));   // src/ram.vhd(56[12:17])
    SB_LUT4 i869_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_28_5), .O(n1117));   // src/ram.vhd(68[19:45])
    defparam i869_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i980_981 (.Q(ram_s_40_2), .C(CLK_3P3_MHZ_c), .D(n1210));   // src/ram.vhd(56[12:17])
    SB_LUT4 i868_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_28_4), .O(n1116));   // src/ram.vhd(68[19:45])
    defparam i868_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i977_978 (.Q(ram_s_40_1), .C(CLK_3P3_MHZ_c), .D(n1209));   // src/ram.vhd(56[12:17])
    SB_LUT4 i867_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_28_3), .O(n1115));   // src/ram.vhd(68[19:45])
    defparam i867_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i974_975 (.Q(ram_s_40_0), .C(CLK_3P3_MHZ_c), .D(n1208));   // src/ram.vhd(56[12:17])
    SB_LUT4 i866_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_28_2), .O(n1114));   // src/ram.vhd(68[19:45])
    defparam i866_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i971_972 (.Q(ram_s_39_7), .C(CLK_3P3_MHZ_c), .D(n1207));   // src/ram.vhd(56[12:17])
    SB_LUT4 i865_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_28_1), .O(n1113));   // src/ram.vhd(68[19:45])
    defparam i865_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i968_969 (.Q(ram_s_39_6), .C(CLK_3P3_MHZ_c), .D(n1206));   // src/ram.vhd(56[12:17])
    SB_LUT4 i864_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_28_0), .O(n1112));   // src/ram.vhd(68[19:45])
    defparam i864_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i965_966 (.Q(ram_s_39_5), .C(CLK_3P3_MHZ_c), .D(n1205));   // src/ram.vhd(56[12:17])
    SB_LUT4 i879_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_29_7), .O(n1127));   // src/ram.vhd(68[19:45])
    defparam i879_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i962_963 (.Q(ram_s_39_4), .C(CLK_3P3_MHZ_c), .D(n1204));   // src/ram.vhd(56[12:17])
    SB_LUT4 i878_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_29_6), .O(n1126));   // src/ram.vhd(68[19:45])
    defparam i878_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i959_960 (.Q(ram_s_39_3), .C(CLK_3P3_MHZ_c), .D(n1203));   // src/ram.vhd(56[12:17])
    SB_LUT4 i877_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_29_5), .O(n1125));   // src/ram.vhd(68[19:45])
    defparam i877_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i956_957 (.Q(ram_s_39_2), .C(CLK_3P3_MHZ_c), .D(n1202));   // src/ram.vhd(56[12:17])
    SB_LUT4 i876_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_29_4), .O(n1124));   // src/ram.vhd(68[19:45])
    defparam i876_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i953_954 (.Q(ram_s_39_1), .C(CLK_3P3_MHZ_c), .D(n1201));   // src/ram.vhd(56[12:17])
    SB_LUT4 i875_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_29_3), .O(n1123));   // src/ram.vhd(68[19:45])
    defparam i875_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i950_951 (.Q(ram_s_39_0), .C(CLK_3P3_MHZ_c), .D(n1200));   // src/ram.vhd(56[12:17])
    SB_LUT4 i874_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_29_2), .O(n1122));   // src/ram.vhd(68[19:45])
    defparam i874_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i947_948 (.Q(ram_s_38_7), .C(CLK_3P3_MHZ_c), .D(n1199));   // src/ram.vhd(56[12:17])
    SB_LUT4 i873_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_29_1), .O(n1121));   // src/ram.vhd(68[19:45])
    defparam i873_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i944_945 (.Q(ram_s_38_6), .C(CLK_3P3_MHZ_c), .D(n1198));   // src/ram.vhd(56[12:17])
    SB_LUT4 i872_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_29_0), .O(n1120));   // src/ram.vhd(68[19:45])
    defparam i872_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i941_942 (.Q(ram_s_38_5), .C(CLK_3P3_MHZ_c), .D(n1197));   // src/ram.vhd(56[12:17])
    SB_LUT4 i887_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_30_7), .O(n1135));   // src/ram.vhd(68[19:45])
    defparam i887_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i938_939 (.Q(ram_s_38_4), .C(CLK_3P3_MHZ_c), .D(n1196));   // src/ram.vhd(56[12:17])
    SB_LUT4 i886_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_30_6), .O(n1134));   // src/ram.vhd(68[19:45])
    defparam i886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i935_936 (.Q(ram_s_38_3), .C(CLK_3P3_MHZ_c), .D(n1195));   // src/ram.vhd(56[12:17])
    SB_LUT4 i885_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_30_5), .O(n1133));   // src/ram.vhd(68[19:45])
    defparam i885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i932_933 (.Q(ram_s_38_2), .C(CLK_3P3_MHZ_c), .D(n1194));   // src/ram.vhd(56[12:17])
    SB_LUT4 i884_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_30_4), .O(n1132));   // src/ram.vhd(68[19:45])
    defparam i884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i929_930 (.Q(ram_s_38_1), .C(CLK_3P3_MHZ_c), .D(n1193));   // src/ram.vhd(56[12:17])
    SB_LUT4 i883_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_30_3), .O(n1131));   // src/ram.vhd(68[19:45])
    defparam i883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i926_927 (.Q(ram_s_38_0), .C(CLK_3P3_MHZ_c), .D(n1192));   // src/ram.vhd(56[12:17])
    SB_LUT4 i882_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_30_2), .O(n1130));   // src/ram.vhd(68[19:45])
    defparam i882_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i923_924 (.Q(ram_s_37_7), .C(CLK_3P3_MHZ_c), .D(n1191));   // src/ram.vhd(56[12:17])
    SB_LUT4 i881_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_30_1), .O(n1129));   // src/ram.vhd(68[19:45])
    defparam i881_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i920_921 (.Q(ram_s_37_6), .C(CLK_3P3_MHZ_c), .D(n1190));   // src/ram.vhd(56[12:17])
    SB_LUT4 i880_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_30_0), .O(n1128));   // src/ram.vhd(68[19:45])
    defparam i880_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i917_918 (.Q(ram_s_37_5), .C(CLK_3P3_MHZ_c), .D(n1189));   // src/ram.vhd(56[12:17])
    SB_LUT4 i895_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_31_7), .O(n1143));   // src/ram.vhd(68[19:45])
    defparam i895_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i914_915 (.Q(ram_s_37_4), .C(CLK_3P3_MHZ_c), .D(n1188));   // src/ram.vhd(56[12:17])
    SB_LUT4 i894_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_31_6), .O(n1142));   // src/ram.vhd(68[19:45])
    defparam i894_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i911_912 (.Q(ram_s_37_3), .C(CLK_3P3_MHZ_c), .D(n1187));   // src/ram.vhd(56[12:17])
    SB_LUT4 i893_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_31_5), .O(n1141));   // src/ram.vhd(68[19:45])
    defparam i893_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i908_909 (.Q(ram_s_37_2), .C(CLK_3P3_MHZ_c), .D(n1186));   // src/ram.vhd(56[12:17])
    SB_LUT4 i892_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_31_4), .O(n1140));   // src/ram.vhd(68[19:45])
    defparam i892_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i905_906 (.Q(ram_s_37_1), .C(CLK_3P3_MHZ_c), .D(n1185));   // src/ram.vhd(56[12:17])
    SB_LUT4 i891_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_31_3), .O(n1139));   // src/ram.vhd(68[19:45])
    defparam i891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i902_903 (.Q(ram_s_37_0), .C(CLK_3P3_MHZ_c), .D(n1184));   // src/ram.vhd(56[12:17])
    SB_LUT4 i890_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_31_2), .O(n1138));   // src/ram.vhd(68[19:45])
    defparam i890_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i899_900 (.Q(ram_s_36_7), .C(CLK_3P3_MHZ_c), .D(n1183));   // src/ram.vhd(56[12:17])
    SB_LUT4 i889_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_31_1), .O(n1137));   // src/ram.vhd(68[19:45])
    defparam i889_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i896_897 (.Q(ram_s_36_6), .C(CLK_3P3_MHZ_c), .D(n1182));   // src/ram.vhd(56[12:17])
    SB_LUT4 i888_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_31_0), .O(n1136));   // src/ram.vhd(68[19:45])
    defparam i888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i893_894 (.Q(ram_s_36_5), .C(CLK_3P3_MHZ_c), .D(n1181));   // src/ram.vhd(56[12:17])
    SB_LUT4 i975_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_41_7), .O(n1223));   // src/ram.vhd(68[19:45])
    defparam i975_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i890_891 (.Q(ram_s_36_4), .C(CLK_3P3_MHZ_c), .D(n1180));   // src/ram.vhd(56[12:17])
    SB_LUT4 i974_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_41_6), .O(n1222));   // src/ram.vhd(68[19:45])
    defparam i974_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i887_888 (.Q(ram_s_36_3), .C(CLK_3P3_MHZ_c), .D(n1179));   // src/ram.vhd(56[12:17])
    SB_LUT4 i973_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_41_5), .O(n1221));   // src/ram.vhd(68[19:45])
    defparam i973_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i884_885 (.Q(ram_s_36_2), .C(CLK_3P3_MHZ_c), .D(n1178));   // src/ram.vhd(56[12:17])
    SB_LUT4 i972_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_41_4), .O(n1220));   // src/ram.vhd(68[19:45])
    defparam i972_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i881_882 (.Q(ram_s_36_1), .C(CLK_3P3_MHZ_c), .D(n1177));   // src/ram.vhd(56[12:17])
    SB_LUT4 i971_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_41_3), .O(n1219));   // src/ram.vhd(68[19:45])
    defparam i971_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i970_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_41_2), .O(n1218));   // src/ram.vhd(68[19:45])
    defparam i970_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i969_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_41_1), .O(n1217));   // src/ram.vhd(68[19:45])
    defparam i969_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i878_879 (.Q(ram_s_36_0), .C(CLK_3P3_MHZ_c), .D(n1176));   // src/ram.vhd(56[12:17])
    SB_DFF i875_876 (.Q(ram_s_35_7), .C(CLK_3P3_MHZ_c), .D(n1175));   // src/ram.vhd(56[12:17])
    SB_LUT4 i968_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_41_0), .O(n1216));   // src/ram.vhd(68[19:45])
    defparam i968_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i872_873 (.Q(ram_s_35_6), .C(CLK_3P3_MHZ_c), .D(n1174));   // src/ram.vhd(56[12:17])
    SB_LUT4 i983_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_42_7), .O(n1231));   // src/ram.vhd(68[19:45])
    defparam i983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i869_870 (.Q(ram_s_35_5), .C(CLK_3P3_MHZ_c), .D(n1173));   // src/ram.vhd(56[12:17])
    SB_LUT4 i982_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_42_6), .O(n1230));   // src/ram.vhd(68[19:45])
    defparam i982_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i866_867 (.Q(ram_s_35_4), .C(CLK_3P3_MHZ_c), .D(n1172));   // src/ram.vhd(56[12:17])
    SB_LUT4 i981_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_42_5), .O(n1229));   // src/ram.vhd(68[19:45])
    defparam i981_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i863_864 (.Q(ram_s_35_3), .C(CLK_3P3_MHZ_c), .D(n1171));   // src/ram.vhd(56[12:17])
    SB_LUT4 i980_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_42_4), .O(n1228));   // src/ram.vhd(68[19:45])
    defparam i980_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i860_861 (.Q(ram_s_35_2), .C(CLK_3P3_MHZ_c), .D(n1170));   // src/ram.vhd(56[12:17])
    SB_LUT4 i979_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_42_3), .O(n1227));   // src/ram.vhd(68[19:45])
    defparam i979_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i857_858 (.Q(ram_s_35_1), .C(CLK_3P3_MHZ_c), .D(n1169));   // src/ram.vhd(56[12:17])
    SB_LUT4 i978_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_42_2), .O(n1226));   // src/ram.vhd(68[19:45])
    defparam i978_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i854_855 (.Q(ram_s_35_0), .C(CLK_3P3_MHZ_c), .D(n1168));   // src/ram.vhd(56[12:17])
    SB_LUT4 i977_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_42_1), .O(n1225));   // src/ram.vhd(68[19:45])
    defparam i977_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i851_852 (.Q(ram_s_34_7), .C(CLK_3P3_MHZ_c), .D(n1167));   // src/ram.vhd(56[12:17])
    SB_LUT4 i976_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_42_0), .O(n1224));   // src/ram.vhd(68[19:45])
    defparam i976_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i848_849 (.Q(ram_s_34_6), .C(CLK_3P3_MHZ_c), .D(n1166));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1015_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_46_7), .O(n1263));   // src/ram.vhd(68[19:45])
    defparam i1015_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i845_846 (.Q(ram_s_34_5), .C(CLK_3P3_MHZ_c), .D(n1165));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1014_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_46_6), .O(n1262));   // src/ram.vhd(68[19:45])
    defparam i1014_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i842_843 (.Q(ram_s_34_4), .C(CLK_3P3_MHZ_c), .D(n1164));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1013_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_46_5), .O(n1261));   // src/ram.vhd(68[19:45])
    defparam i1013_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i839_840 (.Q(ram_s_34_3), .C(CLK_3P3_MHZ_c), .D(n1163));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1012_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_46_4), .O(n1260));   // src/ram.vhd(68[19:45])
    defparam i1012_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i836_837 (.Q(ram_s_34_2), .C(CLK_3P3_MHZ_c), .D(n1162));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1011_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_46_3), .O(n1259));   // src/ram.vhd(68[19:45])
    defparam i1011_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i833_834 (.Q(ram_s_34_1), .C(CLK_3P3_MHZ_c), .D(n1161));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1010_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_46_2), .O(n1258));   // src/ram.vhd(68[19:45])
    defparam i1010_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i830_831 (.Q(ram_s_34_0), .C(CLK_3P3_MHZ_c), .D(n1160));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1009_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_46_1), .O(n1257));   // src/ram.vhd(68[19:45])
    defparam i1009_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i827_828 (.Q(ram_s_33_7), .C(CLK_3P3_MHZ_c), .D(n1159));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1008_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_46_0), .O(n1256));   // src/ram.vhd(68[19:45])
    defparam i1008_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i824_825 (.Q(ram_s_33_6), .C(CLK_3P3_MHZ_c), .D(n1158));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1031_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_48_7), .O(n1279));   // src/ram.vhd(68[19:45])
    defparam i1031_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i821_822 (.Q(ram_s_33_5), .C(CLK_3P3_MHZ_c), .D(n1157));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1030_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_48_6), .O(n1278));   // src/ram.vhd(68[19:45])
    defparam i1030_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i818_819 (.Q(ram_s_33_4), .C(CLK_3P3_MHZ_c), .D(n1156));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1029_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_48_5), .O(n1277));   // src/ram.vhd(68[19:45])
    defparam i1029_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i815_816 (.Q(ram_s_33_3), .C(CLK_3P3_MHZ_c), .D(n1155));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1028_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_48_4), .O(n1276));   // src/ram.vhd(68[19:45])
    defparam i1028_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i812_813 (.Q(ram_s_33_2), .C(CLK_3P3_MHZ_c), .D(n1154));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1027_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_48_3), .O(n1275));   // src/ram.vhd(68[19:45])
    defparam i1027_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i809_810 (.Q(ram_s_33_1), .C(CLK_3P3_MHZ_c), .D(n1153));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1026_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_48_2), .O(n1274));   // src/ram.vhd(68[19:45])
    defparam i1026_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i806_807 (.Q(ram_s_33_0), .C(CLK_3P3_MHZ_c), .D(n1152));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1025_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_48_1), .O(n1273));   // src/ram.vhd(68[19:45])
    defparam i1025_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i803_804 (.Q(ram_s_32_7), .C(CLK_3P3_MHZ_c), .D(n1151));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1024_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_48_0), .O(n1272));   // src/ram.vhd(68[19:45])
    defparam i1024_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i800_801 (.Q(ram_s_32_6), .C(CLK_3P3_MHZ_c), .D(n1150));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1039_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_49_7), .O(n1287));   // src/ram.vhd(68[19:45])
    defparam i1039_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i797_798 (.Q(ram_s_32_5), .C(CLK_3P3_MHZ_c), .D(n1149));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1038_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_49_6), .O(n1286));   // src/ram.vhd(68[19:45])
    defparam i1038_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i794_795 (.Q(ram_s_32_4), .C(CLK_3P3_MHZ_c), .D(n1148));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1037_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_49_5), .O(n1285));   // src/ram.vhd(68[19:45])
    defparam i1037_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i791_792 (.Q(ram_s_32_3), .C(CLK_3P3_MHZ_c), .D(n1147));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1036_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_49_4), .O(n1284));   // src/ram.vhd(68[19:45])
    defparam i1036_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i788_789 (.Q(ram_s_32_2), .C(CLK_3P3_MHZ_c), .D(n1146));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1035_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_49_3), .O(n1283));   // src/ram.vhd(68[19:45])
    defparam i1035_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i785_786 (.Q(ram_s_32_1), .C(CLK_3P3_MHZ_c), .D(n1145));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1034_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_49_2), .O(n1282));   // src/ram.vhd(68[19:45])
    defparam i1034_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i782_783 (.Q(ram_s_32_0), .C(CLK_3P3_MHZ_c), .D(n1144));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1033_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_49_1), .O(n1281));   // src/ram.vhd(68[19:45])
    defparam i1033_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i779_780 (.Q(ram_s_31_7), .C(CLK_3P3_MHZ_c), .D(n1143));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1032_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_49_0), .O(n1280));   // src/ram.vhd(68[19:45])
    defparam i1032_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i776_777 (.Q(ram_s_31_6), .C(CLK_3P3_MHZ_c), .D(n1142));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1047_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_50_7), .O(n1295));   // src/ram.vhd(68[19:45])
    defparam i1047_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i773_774 (.Q(ram_s_31_5), .C(CLK_3P3_MHZ_c), .D(n1141));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1046_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_50_6), .O(n1294));   // src/ram.vhd(68[19:45])
    defparam i1046_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i770_771 (.Q(ram_s_31_4), .C(CLK_3P3_MHZ_c), .D(n1140));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1045_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_50_5), .O(n1293));   // src/ram.vhd(68[19:45])
    defparam i1045_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i767_768 (.Q(ram_s_31_3), .C(CLK_3P3_MHZ_c), .D(n1139));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1044_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_50_4), .O(n1292));   // src/ram.vhd(68[19:45])
    defparam i1044_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i764_765 (.Q(ram_s_31_2), .C(CLK_3P3_MHZ_c), .D(n1138));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1043_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_50_3), .O(n1291));   // src/ram.vhd(68[19:45])
    defparam i1043_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i761_762 (.Q(ram_s_31_1), .C(CLK_3P3_MHZ_c), .D(n1137));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1042_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_50_2), .O(n1290));   // src/ram.vhd(68[19:45])
    defparam i1042_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i758_759 (.Q(ram_s_31_0), .C(CLK_3P3_MHZ_c), .D(n1136));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1041_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_50_1), .O(n1289));   // src/ram.vhd(68[19:45])
    defparam i1041_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i755_756 (.Q(ram_s_30_7), .C(CLK_3P3_MHZ_c), .D(n1135));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1040_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_50_0), .O(n1288));   // src/ram.vhd(68[19:45])
    defparam i1040_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i752_753 (.Q(ram_s_30_6), .C(CLK_3P3_MHZ_c), .D(n1134));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1055_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_51_7), .O(n1303));   // src/ram.vhd(68[19:45])
    defparam i1055_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i749_750 (.Q(ram_s_30_5), .C(CLK_3P3_MHZ_c), .D(n1133));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1054_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_51_6), .O(n1302));   // src/ram.vhd(68[19:45])
    defparam i1054_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i746_747 (.Q(ram_s_30_4), .C(CLK_3P3_MHZ_c), .D(n1132));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1053_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_51_5), .O(n1301));   // src/ram.vhd(68[19:45])
    defparam i1053_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i743_744 (.Q(ram_s_30_3), .C(CLK_3P3_MHZ_c), .D(n1131));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1052_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_51_4), .O(n1300));   // src/ram.vhd(68[19:45])
    defparam i1052_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i740_741 (.Q(ram_s_30_2), .C(CLK_3P3_MHZ_c), .D(n1130));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1051_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_51_3), .O(n1299));   // src/ram.vhd(68[19:45])
    defparam i1051_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i737_738 (.Q(ram_s_30_1), .C(CLK_3P3_MHZ_c), .D(n1129));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1050_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_51_2), .O(n1298));   // src/ram.vhd(68[19:45])
    defparam i1050_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i734_735 (.Q(ram_s_30_0), .C(CLK_3P3_MHZ_c), .D(n1128));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1049_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_51_1), .O(n1297));   // src/ram.vhd(68[19:45])
    defparam i1049_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i731_732 (.Q(ram_s_29_7), .C(CLK_3P3_MHZ_c), .D(n1127));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1048_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_51_0), .O(n1296));   // src/ram.vhd(68[19:45])
    defparam i1048_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i728_729 (.Q(ram_s_29_6), .C(CLK_3P3_MHZ_c), .D(n1126));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1063_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_52_7), .O(n1311));   // src/ram.vhd(68[19:45])
    defparam i1063_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i725_726 (.Q(ram_s_29_5), .C(CLK_3P3_MHZ_c), .D(n1125));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1062_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_52_6), .O(n1310));   // src/ram.vhd(68[19:45])
    defparam i1062_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i722_723 (.Q(ram_s_29_4), .C(CLK_3P3_MHZ_c), .D(n1124));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1061_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_52_5), .O(n1309));   // src/ram.vhd(68[19:45])
    defparam i1061_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i719_720 (.Q(ram_s_29_3), .C(CLK_3P3_MHZ_c), .D(n1123));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1060_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_52_4), .O(n1308));   // src/ram.vhd(68[19:45])
    defparam i1060_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i716_717 (.Q(ram_s_29_2), .C(CLK_3P3_MHZ_c), .D(n1122));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1059_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_52_3), .O(n1307));   // src/ram.vhd(68[19:45])
    defparam i1059_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i713_714 (.Q(ram_s_29_1), .C(CLK_3P3_MHZ_c), .D(n1121));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1058_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_52_2), .O(n1306));   // src/ram.vhd(68[19:45])
    defparam i1058_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i710_711 (.Q(ram_s_29_0), .C(CLK_3P3_MHZ_c), .D(n1120));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1057_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_52_1), .O(n1305));   // src/ram.vhd(68[19:45])
    defparam i1057_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i707_708 (.Q(ram_s_28_7), .C(CLK_3P3_MHZ_c), .D(n1119));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1056_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_52_0), .O(n1304));   // src/ram.vhd(68[19:45])
    defparam i1056_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i704_705 (.Q(ram_s_28_6), .C(CLK_3P3_MHZ_c), .D(n1118));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1071_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_53_7), .O(n1319));   // src/ram.vhd(68[19:45])
    defparam i1071_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i701_702 (.Q(ram_s_28_5), .C(CLK_3P3_MHZ_c), .D(n1117));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1070_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_53_6), .O(n1318));   // src/ram.vhd(68[19:45])
    defparam i1070_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i698_699 (.Q(ram_s_28_4), .C(CLK_3P3_MHZ_c), .D(n1116));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1069_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_53_5), .O(n1317));   // src/ram.vhd(68[19:45])
    defparam i1069_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i695_696 (.Q(ram_s_28_3), .C(CLK_3P3_MHZ_c), .D(n1115));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1068_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_53_4), .O(n1316));   // src/ram.vhd(68[19:45])
    defparam i1068_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i692_693 (.Q(ram_s_28_2), .C(CLK_3P3_MHZ_c), .D(n1114));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1067_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_53_3), .O(n1315));   // src/ram.vhd(68[19:45])
    defparam i1067_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i689_690 (.Q(ram_s_28_1), .C(CLK_3P3_MHZ_c), .D(n1113));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1066_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_53_2), .O(n1314));   // src/ram.vhd(68[19:45])
    defparam i1066_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i686_687 (.Q(ram_s_28_0), .C(CLK_3P3_MHZ_c), .D(n1112));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1065_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_53_1), .O(n1313));   // src/ram.vhd(68[19:45])
    defparam i1065_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i683_684 (.Q(ram_s_27_7), .C(CLK_3P3_MHZ_c), .D(n1111));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1064_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_53_0), .O(n1312));   // src/ram.vhd(68[19:45])
    defparam i1064_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i680_681 (.Q(ram_s_27_6), .C(CLK_3P3_MHZ_c), .D(n1110));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1079_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_54_7), .O(n1327));   // src/ram.vhd(68[19:45])
    defparam i1079_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i677_678 (.Q(ram_s_27_5), .C(CLK_3P3_MHZ_c), .D(n1109));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1078_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_54_6), .O(n1326));   // src/ram.vhd(68[19:45])
    defparam i1078_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i674_675 (.Q(ram_s_27_4), .C(CLK_3P3_MHZ_c), .D(n1108));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1077_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_54_5), .O(n1325));   // src/ram.vhd(68[19:45])
    defparam i1077_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i671_672 (.Q(ram_s_27_3), .C(CLK_3P3_MHZ_c), .D(n1107));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1076_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_54_4), .O(n1324));   // src/ram.vhd(68[19:45])
    defparam i1076_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i668_669 (.Q(ram_s_27_2), .C(CLK_3P3_MHZ_c), .D(n1106));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1075_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_54_3), .O(n1323));   // src/ram.vhd(68[19:45])
    defparam i1075_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i665_666 (.Q(ram_s_27_1), .C(CLK_3P3_MHZ_c), .D(n1105));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1074_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_54_2), .O(n1322));   // src/ram.vhd(68[19:45])
    defparam i1074_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i662_663 (.Q(ram_s_27_0), .C(CLK_3P3_MHZ_c), .D(n1104));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1073_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_54_1), .O(n1321));   // src/ram.vhd(68[19:45])
    defparam i1073_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i659_660 (.Q(ram_s_26_7), .C(CLK_3P3_MHZ_c), .D(n1103));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1072_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_54_0), .O(n1320));   // src/ram.vhd(68[19:45])
    defparam i1072_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i656_657 (.Q(ram_s_26_6), .C(CLK_3P3_MHZ_c), .D(n1102));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1087_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_55_7), .O(n1335));   // src/ram.vhd(68[19:45])
    defparam i1087_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i653_654 (.Q(ram_s_26_5), .C(CLK_3P3_MHZ_c), .D(n1101));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1086_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_55_6), .O(n1334));   // src/ram.vhd(68[19:45])
    defparam i1086_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i650_651 (.Q(ram_s_26_4), .C(CLK_3P3_MHZ_c), .D(n1100));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1085_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_55_5), .O(n1333));   // src/ram.vhd(68[19:45])
    defparam i1085_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i647_648 (.Q(ram_s_26_3), .C(CLK_3P3_MHZ_c), .D(n1099));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1084_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_55_4), .O(n1332));   // src/ram.vhd(68[19:45])
    defparam i1084_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i644_645 (.Q(ram_s_26_2), .C(CLK_3P3_MHZ_c), .D(n1098));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1083_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_55_3), .O(n1331));   // src/ram.vhd(68[19:45])
    defparam i1083_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i641_642 (.Q(ram_s_26_1), .C(CLK_3P3_MHZ_c), .D(n1097));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1082_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_55_2), .O(n1330));   // src/ram.vhd(68[19:45])
    defparam i1082_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i638_639 (.Q(ram_s_26_0), .C(CLK_3P3_MHZ_c), .D(n1096));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1081_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_55_1), .O(n1329));   // src/ram.vhd(68[19:45])
    defparam i1081_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i635_636 (.Q(ram_s_25_7), .C(CLK_3P3_MHZ_c), .D(n1095));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1080_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_55_0), .O(n1328));   // src/ram.vhd(68[19:45])
    defparam i1080_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i632_633 (.Q(ram_s_25_6), .C(CLK_3P3_MHZ_c), .D(n1094));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1095_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_56_7), .O(n1343));   // src/ram.vhd(68[19:45])
    defparam i1095_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i629_630 (.Q(ram_s_25_5), .C(CLK_3P3_MHZ_c), .D(n1093));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1094_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_56_6), .O(n1342));   // src/ram.vhd(68[19:45])
    defparam i1094_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i626_627 (.Q(ram_s_25_4), .C(CLK_3P3_MHZ_c), .D(n1092));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1093_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_56_5), .O(n1341));   // src/ram.vhd(68[19:45])
    defparam i1093_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i623_624 (.Q(ram_s_25_3), .C(CLK_3P3_MHZ_c), .D(n1091));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1092_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_56_4), .O(n1340));   // src/ram.vhd(68[19:45])
    defparam i1092_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i620_621 (.Q(ram_s_25_2), .C(CLK_3P3_MHZ_c), .D(n1090));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1091_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_56_3), .O(n1339));   // src/ram.vhd(68[19:45])
    defparam i1091_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i617_618 (.Q(ram_s_25_1), .C(CLK_3P3_MHZ_c), .D(n1089));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1090_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_56_2), .O(n1338));   // src/ram.vhd(68[19:45])
    defparam i1090_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i614_615 (.Q(ram_s_25_0), .C(CLK_3P3_MHZ_c), .D(n1088));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1089_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_56_1), .O(n1337));   // src/ram.vhd(68[19:45])
    defparam i1089_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i611_612 (.Q(ram_s_24_7), .C(CLK_3P3_MHZ_c), .D(n1087));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1088_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_56_0), .O(n1336));   // src/ram.vhd(68[19:45])
    defparam i1088_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i608_609 (.Q(ram_s_24_6), .C(CLK_3P3_MHZ_c), .D(n1086));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1119_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_59_7), .O(n1367));   // src/ram.vhd(68[19:45])
    defparam i1119_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i605_606 (.Q(ram_s_24_5), .C(CLK_3P3_MHZ_c), .D(n1085));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1118_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_59_6), .O(n1366));   // src/ram.vhd(68[19:45])
    defparam i1118_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i602_603 (.Q(ram_s_24_4), .C(CLK_3P3_MHZ_c), .D(n1084));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1117_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_59_5), .O(n1365));   // src/ram.vhd(68[19:45])
    defparam i1117_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i599_600 (.Q(ram_s_24_3), .C(CLK_3P3_MHZ_c), .D(n1083));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1116_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_59_4), .O(n1364));   // src/ram.vhd(68[19:45])
    defparam i1116_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i596_597 (.Q(ram_s_24_2), .C(CLK_3P3_MHZ_c), .D(n1082));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1115_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_59_3), .O(n1363));   // src/ram.vhd(68[19:45])
    defparam i1115_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i593_594 (.Q(ram_s_24_1), .C(CLK_3P3_MHZ_c), .D(n1081));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1114_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_59_2), .O(n1362));   // src/ram.vhd(68[19:45])
    defparam i1114_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i590_591 (.Q(ram_s_24_0), .C(CLK_3P3_MHZ_c), .D(n1080));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1113_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_59_1), .O(n1361));   // src/ram.vhd(68[19:45])
    defparam i1113_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i587_588 (.Q(ram_s_23_7), .C(CLK_3P3_MHZ_c), .D(n1079));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1112_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_59_0), .O(n1360));   // src/ram.vhd(68[19:45])
    defparam i1112_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i584_585 (.Q(ram_s_23_6), .C(CLK_3P3_MHZ_c), .D(n1078));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1127_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_60_7), .O(n1375));   // src/ram.vhd(68[19:45])
    defparam i1127_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i581_582 (.Q(ram_s_23_5), .C(CLK_3P3_MHZ_c), .D(n1077));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1126_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_60_6), .O(n1374));   // src/ram.vhd(68[19:45])
    defparam i1126_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i578_579 (.Q(ram_s_23_4), .C(CLK_3P3_MHZ_c), .D(n1076));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1125_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_60_5), .O(n1373));   // src/ram.vhd(68[19:45])
    defparam i1125_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i575_576 (.Q(ram_s_23_3), .C(CLK_3P3_MHZ_c), .D(n1075));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1124_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_60_4), .O(n1372));   // src/ram.vhd(68[19:45])
    defparam i1124_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i572_573 (.Q(ram_s_23_2), .C(CLK_3P3_MHZ_c), .D(n1074));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1123_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_60_3), .O(n1371));   // src/ram.vhd(68[19:45])
    defparam i1123_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i569_570 (.Q(ram_s_23_1), .C(CLK_3P3_MHZ_c), .D(n1073));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1122_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_60_2), .O(n1370));   // src/ram.vhd(68[19:45])
    defparam i1122_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i566_567 (.Q(ram_s_23_0), .C(CLK_3P3_MHZ_c), .D(n1072));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1121_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_60_1), .O(n1369));   // src/ram.vhd(68[19:45])
    defparam i1121_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i563_564 (.Q(ram_s_22_7), .C(CLK_3P3_MHZ_c), .D(n1071));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1120_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_60_0), .O(n1368));   // src/ram.vhd(68[19:45])
    defparam i1120_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i560_561 (.Q(ram_s_22_6), .C(CLK_3P3_MHZ_c), .D(n1070));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1135_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_61_7), .O(n1383));   // src/ram.vhd(68[19:45])
    defparam i1135_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i557_558 (.Q(ram_s_22_5), .C(CLK_3P3_MHZ_c), .D(n1069));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1134_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_61_6), .O(n1382));   // src/ram.vhd(68[19:45])
    defparam i1134_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i554_555 (.Q(ram_s_22_4), .C(CLK_3P3_MHZ_c), .D(n1068));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1133_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_61_5), .O(n1381));   // src/ram.vhd(68[19:45])
    defparam i1133_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i551_552 (.Q(ram_s_22_3), .C(CLK_3P3_MHZ_c), .D(n1067));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1132_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_61_4), .O(n1380));   // src/ram.vhd(68[19:45])
    defparam i1132_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i548_549 (.Q(ram_s_22_2), .C(CLK_3P3_MHZ_c), .D(n1066));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1131_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_61_3), .O(n1379));   // src/ram.vhd(68[19:45])
    defparam i1131_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i545_546 (.Q(ram_s_22_1), .C(CLK_3P3_MHZ_c), .D(n1065));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1130_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_61_2), .O(n1378));   // src/ram.vhd(68[19:45])
    defparam i1130_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i542_543 (.Q(ram_s_22_0), .C(CLK_3P3_MHZ_c), .D(n1064));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1129_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_61_1), .O(n1377));   // src/ram.vhd(68[19:45])
    defparam i1129_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i539_540 (.Q(ram_s_21_7), .C(CLK_3P3_MHZ_c), .D(n1063));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1128_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_61_0), .O(n1376));   // src/ram.vhd(68[19:45])
    defparam i1128_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i536_537 (.Q(ram_s_21_6), .C(CLK_3P3_MHZ_c), .D(n1062));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2295_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_206_7), .O(n2543));   // src/ram.vhd(68[19:45])
    defparam i2295_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i533_534 (.Q(ram_s_21_5), .C(CLK_3P3_MHZ_c), .D(n1061));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2294_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_206_6), .O(n2542));   // src/ram.vhd(68[19:45])
    defparam i2294_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i395_396 (.Q(ram_s_15_7), .C(CLK_3P3_MHZ_c), .D(n1060));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2293_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_206_5), .O(n2541));   // src/ram.vhd(68[19:45])
    defparam i2293_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i398_399 (.Q(ram_s_16_0), .C(CLK_3P3_MHZ_c), .D(n1059));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2292_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_206_4), .O(n2540));   // src/ram.vhd(68[19:45])
    defparam i2292_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i401_402 (.Q(ram_s_16_1), .C(CLK_3P3_MHZ_c), .D(n1058));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2291_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_206_3), .O(n2539));   // src/ram.vhd(68[19:45])
    defparam i2291_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i476_477 (.Q(ram_s_19_2), .C(CLK_3P3_MHZ_c), .D(n1057));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2290_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_206_2), .O(n2538));   // src/ram.vhd(68[19:45])
    defparam i2290_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i530_531 (.Q(ram_s_21_4), .C(CLK_3P3_MHZ_c), .D(n1056));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2289_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_206_1), .O(n2537));   // src/ram.vhd(68[19:45])
    defparam i2289_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i404_405 (.Q(ram_s_16_2), .C(CLK_3P3_MHZ_c), .D(n1055));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2288_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_206_0), .O(n2536));   // src/ram.vhd(68[19:45])
    defparam i2288_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i407_408 (.Q(ram_s_16_3), .C(CLK_3P3_MHZ_c), .D(n1054));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2287_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_205_7), .O(n2535));   // src/ram.vhd(68[19:45])
    defparam i2287_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i410_411 (.Q(ram_s_16_4), .C(CLK_3P3_MHZ_c), .D(n1053));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2286_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_205_6), .O(n2534));   // src/ram.vhd(68[19:45])
    defparam i2286_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i389_390 (.Q(ram_s_15_5), .C(CLK_3P3_MHZ_c), .D(n1052));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2285_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_205_5), .O(n2533));   // src/ram.vhd(68[19:45])
    defparam i2285_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i365_366 (.Q(ram_s_14_5), .C(CLK_3P3_MHZ_c), .D(n1051));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2284_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_205_4), .O(n2532));   // src/ram.vhd(68[19:45])
    defparam i2284_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i479_480 (.Q(ram_s_19_3), .C(CLK_3P3_MHZ_c), .D(n1050));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2283_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_205_3), .O(n2531));   // src/ram.vhd(68[19:45])
    defparam i2283_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i392_393 (.Q(ram_s_15_6), .C(CLK_3P3_MHZ_c), .D(n1049));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2282_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_205_2), .O(n2530));   // src/ram.vhd(68[19:45])
    defparam i2282_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i413_414 (.Q(ram_s_16_5), .C(CLK_3P3_MHZ_c), .D(n1048));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2281_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_205_1), .O(n2529));   // src/ram.vhd(68[19:45])
    defparam i2281_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i14_15 (.Q(ram_s_0_0), .C(CLK_3P3_MHZ_c), .D(n1047));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2280_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_205_0), .O(n2528));   // src/ram.vhd(68[19:45])
    defparam i2280_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i17_18 (.Q(ram_s_0_1), .C(CLK_3P3_MHZ_c), .D(n1046));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2279_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_204_7), .O(n2527));   // src/ram.vhd(68[19:45])
    defparam i2279_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i20_21 (.Q(ram_s_0_2), .C(CLK_3P3_MHZ_c), .D(n1045));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2278_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_204_6), .O(n2526));   // src/ram.vhd(68[19:45])
    defparam i2278_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i311_312 (.Q(ram_s_12_3), .C(CLK_3P3_MHZ_c), .D(n1044));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2277_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_204_5), .O(n2525));   // src/ram.vhd(68[19:45])
    defparam i2277_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i296_297 (.Q(ram_s_11_6), .C(CLK_3P3_MHZ_c), .D(n1043));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2276_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_204_4), .O(n2524));   // src/ram.vhd(68[19:45])
    defparam i2276_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i281_282 (.Q(ram_s_11_1), .C(CLK_3P3_MHZ_c), .D(n1042));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2275_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_204_3), .O(n2523));   // src/ram.vhd(68[19:45])
    defparam i2275_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i320_321 (.Q(ram_s_12_6), .C(CLK_3P3_MHZ_c), .D(n1041));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2274_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_204_2), .O(n2522));   // src/ram.vhd(68[19:45])
    defparam i2274_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i305_306 (.Q(ram_s_12_1), .C(CLK_3P3_MHZ_c), .D(n1040));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2273_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_204_1), .O(n2521));   // src/ram.vhd(68[19:45])
    defparam i2273_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i440_441 (.Q(ram_s_17_6), .C(CLK_3P3_MHZ_c), .D(n1039));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2272_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_204_0), .O(n2520));   // src/ram.vhd(68[19:45])
    defparam i2272_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i290_291 (.Q(ram_s_11_4), .C(CLK_3P3_MHZ_c), .D(n1038));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i414_2_lut_3_lut (.I0(n94_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n182));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i414_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i314_315 (.Q(ram_s_12_4), .C(CLK_3P3_MHZ_c), .D(n1037));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i413_2_lut_3_lut (.I0(n94_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n54));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i413_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i299_300 (.Q(ram_s_11_7), .C(CLK_3P3_MHZ_c), .D(n1036));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i412_2_lut_3_lut (.I0(n92_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n183));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i412_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i284_285 (.Q(ram_s_11_2), .C(CLK_3P3_MHZ_c), .D(n1035));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i411_2_lut_3_lut (.I0(n92_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n55));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i411_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i323_324 (.Q(ram_s_12_7), .C(CLK_3P3_MHZ_c), .D(n1034));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i410_2_lut_3_lut (.I0(n90_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n184));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i410_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i308_309 (.Q(ram_s_12_2), .C(CLK_3P3_MHZ_c), .D(n1033));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i409_2_lut_3_lut (.I0(n90_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n56));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i409_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i293_294 (.Q(ram_s_11_5), .C(CLK_3P3_MHZ_c), .D(n1032));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i408_2_lut_3_lut (.I0(n88), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n185));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i408_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i317_318 (.Q(ram_s_12_5), .C(CLK_3P3_MHZ_c), .D(n1031));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i407_2_lut_3_lut (.I0(n88), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n57));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i407_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i302_303 (.Q(ram_s_12_0), .C(CLK_3P3_MHZ_c), .D(n1030));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i406_2_lut_3_lut (.I0(n86_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n186));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i406_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i287_288 (.Q(ram_s_11_3), .C(CLK_3P3_MHZ_c), .D(n1029));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i405_2_lut_3_lut (.I0(n86_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n58));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i405_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i482_483 (.Q(ram_s_19_4), .C(CLK_3P3_MHZ_c), .D(n1028));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i404_2_lut_3_lut (.I0(n84_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n187));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i404_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i485_486 (.Q(ram_s_19_5), .C(CLK_3P3_MHZ_c), .D(n1027));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i403_2_lut_3_lut (.I0(n84_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n59));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i403_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i488_489 (.Q(ram_s_19_6), .C(CLK_3P3_MHZ_c), .D(n1026));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i402_2_lut_3_lut (.I0(n82_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n188));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i402_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i491_492 (.Q(ram_s_19_7), .C(CLK_3P3_MHZ_c), .D(n1025));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i401_2_lut_3_lut (.I0(n82_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n60));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i401_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i452_453 (.Q(ram_s_18_2), .C(CLK_3P3_MHZ_c), .D(n1024));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i400_2_lut_3_lut (.I0(n80), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n189));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i400_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i455_456 (.Q(ram_s_18_3), .C(CLK_3P3_MHZ_c), .D(n1023));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i399_2_lut_3_lut (.I0(n80), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n61));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i399_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i458_459 (.Q(ram_s_18_4), .C(CLK_3P3_MHZ_c), .D(n1022));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i398_2_lut_3_lut (.I0(n78), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n190));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i398_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i461_462 (.Q(ram_s_18_5), .C(CLK_3P3_MHZ_c), .D(n1021));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i397_2_lut_3_lut (.I0(n78), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n62));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i397_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i464_465 (.Q(ram_s_18_6), .C(CLK_3P3_MHZ_c), .D(n1020));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i396_2_lut_3_lut (.I0(n76), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n191));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i396_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i467_468 (.Q(ram_s_18_7), .C(CLK_3P3_MHZ_c), .D(n1019));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i395_2_lut_3_lut (.I0(n76), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n63));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i395_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i470_471 (.Q(ram_s_19_0), .C(CLK_3P3_MHZ_c), .D(n1018));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i394_2_lut_3_lut (.I0(n74), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n192));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i394_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i23_24 (.Q(ram_s_0_3), .C(CLK_3P3_MHZ_c), .D(n1017));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i393_2_lut_3_lut (.I0(n74), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n64));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i393_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i26_27 (.Q(ram_s_0_4), .C(CLK_3P3_MHZ_c), .D(n1016));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i392_2_lut_3_lut (.I0(n72_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n193));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i392_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i29_30 (.Q(ram_s_0_5), .C(CLK_3P3_MHZ_c), .D(n1015));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i391_2_lut_3_lut (.I0(n72_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n65));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i391_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i32_33 (.Q(ram_s_0_6), .C(CLK_3P3_MHZ_c), .D(n1014));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i390_2_lut_3_lut (.I0(n133), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n194));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i390_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i35_36 (.Q(ram_s_0_7), .C(CLK_3P3_MHZ_c), .D(n1013));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i389_2_lut_3_lut (.I0(n133), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n66));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i389_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i38_39 (.Q(ram_s_1_0), .C(CLK_3P3_MHZ_c), .D(n1012));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i388_2_lut_3_lut (.I0(n131), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n195));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i388_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i41_42 (.Q(ram_s_1_1), .C(CLK_3P3_MHZ_c), .D(n1011));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i387_2_lut_3_lut (.I0(n131), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n67));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i387_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i44_45 (.Q(ram_s_1_2), .C(CLK_3P3_MHZ_c), .D(n1010));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2159_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_189_7), .O(n2407));   // src/ram.vhd(68[19:45])
    defparam i2159_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i47_48 (.Q(ram_s_1_3), .C(CLK_3P3_MHZ_c), .D(n1009));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2158_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_189_6), .O(n2406));   // src/ram.vhd(68[19:45])
    defparam i2158_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i50_51 (.Q(ram_s_1_4), .C(CLK_3P3_MHZ_c), .D(n1008));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2157_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_189_5), .O(n2405));   // src/ram.vhd(68[19:45])
    defparam i2157_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i53_54 (.Q(ram_s_1_5), .C(CLK_3P3_MHZ_c), .D(n1007));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2156_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_189_4), .O(n2404));   // src/ram.vhd(68[19:45])
    defparam i2156_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i122_123 (.Q(ram_s_4_4), .C(CLK_3P3_MHZ_c), .D(n1006));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2155_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_189_3), .O(n2403));   // src/ram.vhd(68[19:45])
    defparam i2155_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i131_132 (.Q(ram_s_4_7), .C(CLK_3P3_MHZ_c), .D(n1005));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2154_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_189_2), .O(n2402));   // src/ram.vhd(68[19:45])
    defparam i2154_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i125_126 (.Q(ram_s_4_5), .C(CLK_3P3_MHZ_c), .D(n1004));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2153_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_189_1), .O(n2401));   // src/ram.vhd(68[19:45])
    defparam i2153_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i134_135 (.Q(ram_s_5_0), .C(CLK_3P3_MHZ_c), .D(n1003));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2152_3_lut_4_lut (.I0(n258), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_189_0), .O(n2400));   // src/ram.vhd(68[19:45])
    defparam i2152_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i128_129 (.Q(ram_s_4_6), .C(CLK_3P3_MHZ_c), .D(n1002));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2151_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_188_7), .O(n2399));   // src/ram.vhd(68[19:45])
    defparam i2151_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i137_138 (.Q(ram_s_5_1), .C(CLK_3P3_MHZ_c), .D(n1001));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2150_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_188_6), .O(n2398));   // src/ram.vhd(68[19:45])
    defparam i2150_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i239_240 (.Q(ram_s_9_3), .C(CLK_3P3_MHZ_c), .D(n1000));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2149_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_188_5), .O(n2397));   // src/ram.vhd(68[19:45])
    defparam i2149_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i230_231 (.Q(ram_s_9_0), .C(CLK_3P3_MHZ_c), .D(n999));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2148_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_188_4), .O(n2396));   // src/ram.vhd(68[19:45])
    defparam i2148_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i221_222 (.Q(ram_s_8_5), .C(CLK_3P3_MHZ_c), .D(n998));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2147_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_188_3), .O(n2395));   // src/ram.vhd(68[19:45])
    defparam i2147_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i212_213 (.Q(ram_s_8_2), .C(CLK_3P3_MHZ_c), .D(n997));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2146_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_188_2), .O(n2394));   // src/ram.vhd(68[19:45])
    defparam i2146_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i203_204 (.Q(ram_s_7_7), .C(CLK_3P3_MHZ_c), .D(n996));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2145_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_188_1), .O(n2393));   // src/ram.vhd(68[19:45])
    defparam i2145_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i194_195 (.Q(ram_s_7_4), .C(CLK_3P3_MHZ_c), .D(n995));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2144_3_lut_4_lut (.I0(n256_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_188_0), .O(n2392));   // src/ram.vhd(68[19:45])
    defparam i2144_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i185_186 (.Q(ram_s_7_1), .C(CLK_3P3_MHZ_c), .D(n994));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2143_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_187_7), .O(n2391));   // src/ram.vhd(68[19:45])
    defparam i2143_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i176_177 (.Q(ram_s_6_6), .C(CLK_3P3_MHZ_c), .D(n993));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2142_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_187_6), .O(n2390));   // src/ram.vhd(68[19:45])
    defparam i2142_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i167_168 (.Q(ram_s_6_3), .C(CLK_3P3_MHZ_c), .D(n992));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2141_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_187_5), .O(n2389));   // src/ram.vhd(68[19:45])
    defparam i2141_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i242_243 (.Q(ram_s_9_4), .C(CLK_3P3_MHZ_c), .D(n991));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2140_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_187_4), .O(n2388));   // src/ram.vhd(68[19:45])
    defparam i2140_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i233_234 (.Q(ram_s_9_1), .C(CLK_3P3_MHZ_c), .D(n990));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2139_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_187_3), .O(n2387));   // src/ram.vhd(68[19:45])
    defparam i2139_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i224_225 (.Q(ram_s_8_6), .C(CLK_3P3_MHZ_c), .D(n989));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2138_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_187_2), .O(n2386));   // src/ram.vhd(68[19:45])
    defparam i2138_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i215_216 (.Q(ram_s_8_3), .C(CLK_3P3_MHZ_c), .D(n988));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2137_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_187_1), .O(n2385));   // src/ram.vhd(68[19:45])
    defparam i2137_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i206_207 (.Q(ram_s_8_0), .C(CLK_3P3_MHZ_c), .D(n987));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2136_3_lut_4_lut (.I0(n254_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_187_0), .O(n2384));   // src/ram.vhd(68[19:45])
    defparam i2136_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i197_198 (.Q(ram_s_7_5), .C(CLK_3P3_MHZ_c), .D(n986));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i380_2_lut_3_lut (.I0(n123_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n199));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i380_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i188_189 (.Q(ram_s_7_2), .C(CLK_3P3_MHZ_c), .D(n985));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i379_2_lut_3_lut (.I0(n123_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n71));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i379_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i179_180 (.Q(ram_s_6_7), .C(CLK_3P3_MHZ_c), .D(n984));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i378_2_lut_3_lut (.I0(n121_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n200));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i378_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i170_171 (.Q(ram_s_6_4), .C(CLK_3P3_MHZ_c), .D(n983));   // src/ram.vhd(56[12:17])
    SB_LUT4 EnabledDecoder_2_i377_2_lut_3_lut (.I0(n121_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n72));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i377_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i245_246 (.Q(ram_s_9_5), .C(CLK_3P3_MHZ_c), .D(n982));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2119_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_184_7), .O(n2367));   // src/ram.vhd(68[19:45])
    defparam i2119_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i236_237 (.Q(ram_s_9_2), .C(CLK_3P3_MHZ_c), .D(n981));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2118_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_184_6), .O(n2366));   // src/ram.vhd(68[19:45])
    defparam i2118_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i227_228 (.Q(ram_s_8_7), .C(CLK_3P3_MHZ_c), .D(n980));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2117_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_184_5), .O(n2365));   // src/ram.vhd(68[19:45])
    defparam i2117_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i218_219 (.Q(ram_s_8_4), .C(CLK_3P3_MHZ_c), .D(n979));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2116_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_184_4), .O(n2364));   // src/ram.vhd(68[19:45])
    defparam i2116_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i209_210 (.Q(ram_s_8_1), .C(CLK_3P3_MHZ_c), .D(n978));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2115_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_184_3), .O(n2363));   // src/ram.vhd(68[19:45])
    defparam i2115_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i200_201 (.Q(ram_s_7_6), .C(CLK_3P3_MHZ_c), .D(n977));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2114_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_184_2), .O(n2362));   // src/ram.vhd(68[19:45])
    defparam i2114_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i191_192 (.Q(ram_s_7_3), .C(CLK_3P3_MHZ_c), .D(n976));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2113_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_184_1), .O(n2361));   // src/ram.vhd(68[19:45])
    defparam i2113_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i182_183 (.Q(ram_s_7_0), .C(CLK_3P3_MHZ_c), .D(n975));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2112_3_lut_4_lut (.I0(n248), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_184_0), .O(n2360));   // src/ram.vhd(68[19:45])
    defparam i2112_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i173_174 (.Q(ram_s_6_5), .C(CLK_3P3_MHZ_c), .D(n974));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2111_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_183_7), .O(n2359));   // src/ram.vhd(68[19:45])
    defparam i2111_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i56_57 (.Q(ram_s_1_6), .C(CLK_3P3_MHZ_c), .D(n973));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2110_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_183_6), .O(n2358));   // src/ram.vhd(68[19:45])
    defparam i2110_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i59_60 (.Q(ram_s_1_7), .C(CLK_3P3_MHZ_c), .D(n972));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2109_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_183_5), .O(n2357));   // src/ram.vhd(68[19:45])
    defparam i2109_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i62_63 (.Q(ram_s_2_0), .C(CLK_3P3_MHZ_c), .D(n971));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2108_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_183_4), .O(n2356));   // src/ram.vhd(68[19:45])
    defparam i2108_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i65_66 (.Q(ram_s_2_1), .C(CLK_3P3_MHZ_c), .D(n970));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2107_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_183_3), .O(n2355));   // src/ram.vhd(68[19:45])
    defparam i2107_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i68_69 (.Q(ram_s_2_2), .C(CLK_3P3_MHZ_c), .D(n969));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2106_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_183_2), .O(n2354));   // src/ram.vhd(68[19:45])
    defparam i2106_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i71_72 (.Q(ram_s_2_3), .C(CLK_3P3_MHZ_c), .D(n968));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2105_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_183_1), .O(n2353));   // src/ram.vhd(68[19:45])
    defparam i2105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i74_75 (.Q(ram_s_2_4), .C(CLK_3P3_MHZ_c), .D(n967));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2104_3_lut_4_lut (.I0(n246_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_183_0), .O(n2352));   // src/ram.vhd(68[19:45])
    defparam i2104_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i77_78 (.Q(ram_s_2_5), .C(CLK_3P3_MHZ_c), .D(n966));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2103_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_182_7), .O(n2351));   // src/ram.vhd(68[19:45])
    defparam i2103_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i80_81 (.Q(ram_s_2_6), .C(CLK_3P3_MHZ_c), .D(n965));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2102_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_182_6), .O(n2350));   // src/ram.vhd(68[19:45])
    defparam i2102_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i83_84 (.Q(ram_s_2_7), .C(CLK_3P3_MHZ_c), .D(n964));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2101_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_182_5), .O(n2349));   // src/ram.vhd(68[19:45])
    defparam i2101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i86_87 (.Q(ram_s_3_0), .C(CLK_3P3_MHZ_c), .D(n963));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2100_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_182_4), .O(n2348));   // src/ram.vhd(68[19:45])
    defparam i2100_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i89_90 (.Q(ram_s_3_1), .C(CLK_3P3_MHZ_c), .D(n962));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2099_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_182_3), .O(n2347));   // src/ram.vhd(68[19:45])
    defparam i2099_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i92_93 (.Q(ram_s_3_2), .C(CLK_3P3_MHZ_c), .D(n961));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2098_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_182_2), .O(n2346));   // src/ram.vhd(68[19:45])
    defparam i2098_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i95_96 (.Q(ram_s_3_3), .C(CLK_3P3_MHZ_c), .D(n960));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2097_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_182_1), .O(n2345));   // src/ram.vhd(68[19:45])
    defparam i2097_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i98_99 (.Q(ram_s_3_4), .C(CLK_3P3_MHZ_c), .D(n959));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2096_3_lut_4_lut (.I0(n244_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_182_0), .O(n2344));   // src/ram.vhd(68[19:45])
    defparam i2096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i101_102 (.Q(ram_s_3_5), .C(CLK_3P3_MHZ_c), .D(n958));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2095_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_181_7), .O(n2343));   // src/ram.vhd(68[19:45])
    defparam i2095_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i371_372 (.Q(ram_s_14_7), .C(CLK_3P3_MHZ_c), .D(n957));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2094_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_181_6), .O(n2342));   // src/ram.vhd(68[19:45])
    defparam i2094_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i374_375 (.Q(ram_s_15_0), .C(CLK_3P3_MHZ_c), .D(n956));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2093_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_181_5), .O(n2341));   // src/ram.vhd(68[19:45])
    defparam i2093_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i494_495 (.Q(ram_s_20_0), .C(CLK_3P3_MHZ_c), .D(n955));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2092_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_181_4), .O(n2340));   // src/ram.vhd(68[19:45])
    defparam i2092_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i497_498 (.Q(ram_s_20_1), .C(CLK_3P3_MHZ_c), .D(n954));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2091_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_181_3), .O(n2339));   // src/ram.vhd(68[19:45])
    defparam i2091_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i416_417 (.Q(ram_s_16_6), .C(CLK_3P3_MHZ_c), .D(n953));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2090_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_181_2), .O(n2338));   // src/ram.vhd(68[19:45])
    defparam i2090_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i104_105 (.Q(ram_s_3_6), .C(CLK_3P3_MHZ_c), .D(n952));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2089_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_181_1), .O(n2337));   // src/ram.vhd(68[19:45])
    defparam i2089_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i419_420 (.Q(ram_s_16_7), .C(CLK_3P3_MHZ_c), .D(n951));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2088_3_lut_4_lut (.I0(n242), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_181_0), .O(n2336));   // src/ram.vhd(68[19:45])
    defparam i2088_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i107_108 (.Q(ram_s_3_7), .C(CLK_3P3_MHZ_c), .D(n950));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2087_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_180_7), .O(n2335));   // src/ram.vhd(68[19:45])
    defparam i2087_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i269_270 (.Q(ram_s_10_5), .C(CLK_3P3_MHZ_c), .D(n949));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2086_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_180_6), .O(n2334));   // src/ram.vhd(68[19:45])
    defparam i2086_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i272_273 (.Q(ram_s_10_6), .C(CLK_3P3_MHZ_c), .D(n948));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2085_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_180_5), .O(n2333));   // src/ram.vhd(68[19:45])
    defparam i2085_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i500_501 (.Q(ram_s_20_2), .C(CLK_3P3_MHZ_c), .D(n947));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2084_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_180_4), .O(n2332));   // src/ram.vhd(68[19:45])
    defparam i2084_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i110_111 (.Q(ram_s_4_0), .C(CLK_3P3_MHZ_c), .D(n946));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2083_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_180_3), .O(n2331));   // src/ram.vhd(68[19:45])
    defparam i2083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i503_504 (.Q(ram_s_20_3), .C(CLK_3P3_MHZ_c), .D(n945));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2082_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_180_2), .O(n2330));   // src/ram.vhd(68[19:45])
    defparam i2082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i113_114 (.Q(ram_s_4_1), .C(CLK_3P3_MHZ_c), .D(n944));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2081_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_180_1), .O(n2329));   // src/ram.vhd(68[19:45])
    defparam i2081_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i506_507 (.Q(ram_s_20_4), .C(CLK_3P3_MHZ_c), .D(n943));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2080_3_lut_4_lut (.I0(n240), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_180_0), .O(n2328));   // src/ram.vhd(68[19:45])
    defparam i2080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i509_510 (.Q(ram_s_20_5), .C(CLK_3P3_MHZ_c), .D(n942));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2079_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_179_7), .O(n2327));   // src/ram.vhd(68[19:45])
    defparam i2079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i116_117 (.Q(ram_s_4_2), .C(CLK_3P3_MHZ_c), .D(n941));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2078_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_179_6), .O(n2326));   // src/ram.vhd(68[19:45])
    defparam i2078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i140_141 (.Q(ram_s_5_2), .C(CLK_3P3_MHZ_c), .D(n940));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2077_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_179_5), .O(n2325));   // src/ram.vhd(68[19:45])
    defparam i2077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i143_144 (.Q(ram_s_5_3), .C(CLK_3P3_MHZ_c), .D(n939));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2076_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_179_4), .O(n2324));   // src/ram.vhd(68[19:45])
    defparam i2076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i149_150 (.Q(ram_s_5_5), .C(CLK_3P3_MHZ_c), .D(n935));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2075_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_179_3), .O(n2323));   // src/ram.vhd(68[19:45])
    defparam i2075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2074_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_179_2), .O(n2322));   // src/ram.vhd(68[19:45])
    defparam i2074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2073_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_179_1), .O(n2321));   // src/ram.vhd(68[19:45])
    defparam i2073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2072_3_lut_4_lut (.I0(n238), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_179_0), .O(n2320));   // src/ram.vhd(68[19:45])
    defparam i2072_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2071_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_178_7), .O(n2319));   // src/ram.vhd(68[19:45])
    defparam i2071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2322_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_210_2), .O(n2570));   // src/ram.vhd(68[19:45])
    defparam i2322_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2070_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_178_6), .O(n2318));   // src/ram.vhd(68[19:45])
    defparam i2070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i158_159 (.Q(ram_s_6_0), .C(CLK_3P3_MHZ_c), .D(n934));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2069_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_178_5), .O(n2317));   // src/ram.vhd(68[19:45])
    defparam i2069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i161_162 (.Q(ram_s_6_1), .C(CLK_3P3_MHZ_c), .D(n933));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2068_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_178_4), .O(n2316));   // src/ram.vhd(68[19:45])
    defparam i2068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i164_165 (.Q(ram_s_6_2), .C(CLK_3P3_MHZ_c), .D(n932));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2067_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_178_3), .O(n2315));   // src/ram.vhd(68[19:45])
    defparam i2067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i152_153 (.Q(ram_s_5_6), .C(CLK_3P3_MHZ_c), .D(n931));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2066_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_178_2), .O(n2314));   // src/ram.vhd(68[19:45])
    defparam i2066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i155_156 (.Q(ram_s_5_7), .C(CLK_3P3_MHZ_c), .D(n930));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2065_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_178_1), .O(n2313));   // src/ram.vhd(68[19:45])
    defparam i2065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i512_513 (.Q(ram_s_20_6), .C(CLK_3P3_MHZ_c), .D(n929));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2064_3_lut_4_lut (.I0(n236), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_178_0), .O(n2312));   // src/ram.vhd(68[19:45])
    defparam i2064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i251_252 (.Q(ram_s_9_7), .C(CLK_3P3_MHZ_c), .D(n928));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2063_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_177_7), .O(n2311));   // src/ram.vhd(68[19:45])
    defparam i2063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i119_120 (.Q(ram_s_4_3), .C(CLK_3P3_MHZ_c), .D(n927));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2062_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_177_6), .O(n2310));   // src/ram.vhd(68[19:45])
    defparam i2062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i341_342 (.Q(ram_s_13_5), .C(CLK_3P3_MHZ_c), .D(n926));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2061_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_177_5), .O(n2309));   // src/ram.vhd(68[19:45])
    defparam i2061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i335_336 (.Q(ram_s_13_3), .C(CLK_3P3_MHZ_c), .D(n925));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2060_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_177_4), .O(n2308));   // src/ram.vhd(68[19:45])
    defparam i2060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i338_339 (.Q(ram_s_13_4), .C(CLK_3P3_MHZ_c), .D(n924));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2059_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_177_3), .O(n2307));   // src/ram.vhd(68[19:45])
    defparam i2059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i344_345 (.Q(ram_s_13_6), .C(CLK_3P3_MHZ_c), .D(n923));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2058_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_177_2), .O(n2306));   // src/ram.vhd(68[19:45])
    defparam i2058_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i515_516 (.Q(ram_s_20_7), .C(CLK_3P3_MHZ_c), .D(n922));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2057_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_177_1), .O(n2305));   // src/ram.vhd(68[19:45])
    defparam i2057_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2056_3_lut_4_lut (.I0(n234), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_177_0), .O(n2304));   // src/ram.vhd(68[19:45])
    defparam i2056_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2055_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_176_7), .O(n2303));   // src/ram.vhd(68[19:45])
    defparam i2055_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2054_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_176_6), .O(n2302));   // src/ram.vhd(68[19:45])
    defparam i2054_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2491_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_231_3), .O(n2739));   // src/ram.vhd(68[19:45])
    defparam i2491_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2053_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_176_5), .O(n2301));   // src/ram.vhd(68[19:45])
    defparam i2053_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2052_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_176_4), .O(n2300));   // src/ram.vhd(68[19:45])
    defparam i2052_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2051_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_176_3), .O(n2299));   // src/ram.vhd(68[19:45])
    defparam i2051_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2050_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_176_2), .O(n2298));   // src/ram.vhd(68[19:45])
    defparam i2050_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2049_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_176_1), .O(n2297));   // src/ram.vhd(68[19:45])
    defparam i2049_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2048_3_lut_4_lut (.I0(n232), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_176_0), .O(n2296));   // src/ram.vhd(68[19:45])
    defparam i2048_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i358_2_lut_3_lut (.I0(n101), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n210));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i358_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i357_2_lut_3_lut (.I0(n101), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n82));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i357_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2490_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_231_2), .O(n2738));   // src/ram.vhd(68[19:45])
    defparam i2490_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2489_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_231_1), .O(n2737));   // src/ram.vhd(68[19:45])
    defparam i2489_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2488_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_231_0), .O(n2736));   // src/ram.vhd(68[19:45])
    defparam i2488_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2039_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_174_7), .O(n2287));   // src/ram.vhd(68[19:45])
    defparam i2039_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2038_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_174_6), .O(n2286));   // src/ram.vhd(68[19:45])
    defparam i2038_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2037_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_174_5), .O(n2285));   // src/ram.vhd(68[19:45])
    defparam i2037_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2036_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_174_4), .O(n2284));   // src/ram.vhd(68[19:45])
    defparam i2036_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2035_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_174_3), .O(n2283));   // src/ram.vhd(68[19:45])
    defparam i2035_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2034_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_174_2), .O(n2282));   // src/ram.vhd(68[19:45])
    defparam i2034_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2033_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_174_1), .O(n2281));   // src/ram.vhd(68[19:45])
    defparam i2033_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_1__bdd_4_lut_10392 (.I0(port_id[1]), .I1(n9375), .I2(n9376), 
            .I3(port_id[2]), .O(n11465));
    defparam port_id_1__bdd_4_lut_10392.LUT_INIT = 16'he4aa;
    SB_LUT4 n11465_bdd_4_lut (.I0(n11465), .I1(n9352), .I2(n9351), .I3(port_id[2]), 
            .O(n11468));
    defparam n11465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut_10611 (.I0(port_id[3]), .I1(n10104), .I2(n10105), 
            .I3(port_id[4]), .O(n11459));
    defparam port_id_3__bdd_4_lut_10611.LUT_INIT = 16'he4aa;
    SB_LUT4 n11459_bdd_4_lut (.I0(n11459), .I1(n10102), .I2(n10101), .I3(port_id[4]), 
            .O(n11462));
    defparam n11459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10362 (.I0(port_id[0]), .I1(ram_s_42_0), 
            .I2(ram_s_43_0), .I3(port_id[1]), .O(n11453));
    defparam port_id_0__bdd_4_lut_10362.LUT_INIT = 16'he4aa;
    SB_LUT4 n11453_bdd_4_lut (.I0(n11453), .I1(ram_s_41_0), .I2(ram_s_40_0), 
            .I3(port_id[1]), .O(n11456));
    defparam n11453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_10352 (.I0(port_id[1]), .I1(n9306), .I2(n9307), 
            .I3(port_id[2]), .O(n11447));
    defparam port_id_1__bdd_4_lut_10352.LUT_INIT = 16'he4aa;
    SB_LUT4 n11447_bdd_4_lut (.I0(n11447), .I1(n9292), .I2(n9291), .I3(port_id[2]), 
            .O(n11450));
    defparam n11447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10412 (.I0(port_id[2]), .I1(n10439), .I2(n10475), 
            .I3(port_id[3]), .O(n11441));
    defparam port_id_2__bdd_4_lut_10412.LUT_INIT = 16'he4aa;
    SB_LUT4 n11441_bdd_4_lut (.I0(n11441), .I1(n10418), .I2(n10388), .I3(port_id[3]), 
            .O(n11444));
    defparam n11441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10343 (.I0(port_id[0]), .I1(ram_s_198_1), 
            .I2(ram_s_199_1), .I3(port_id[1]), .O(n11429));
    defparam port_id_0__bdd_4_lut_10343.LUT_INIT = 16'he4aa;
    SB_LUT4 n11429_bdd_4_lut (.I0(n11429), .I1(ram_s_197_1), .I2(ram_s_196_1), 
            .I3(port_id[1]), .O(n11432));
    defparam n11429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10323 (.I0(port_id[0]), .I1(ram_s_194_2), 
            .I2(ram_s_195_2), .I3(port_id[1]), .O(n11423));
    defparam port_id_0__bdd_4_lut_10323.LUT_INIT = 16'he4aa;
    SB_LUT4 n11423_bdd_4_lut (.I0(n11423), .I1(ram_s_193_2), .I2(ram_s_192_2), 
            .I3(port_id[1]), .O(n11426));
    defparam n11423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10333 (.I0(port_id[2]), .I1(n10613), .I2(n10631), 
            .I3(port_id[3]), .O(n11417));
    defparam port_id_2__bdd_4_lut_10333.LUT_INIT = 16'he4aa;
    SB_LUT4 n11417_bdd_4_lut (.I0(n11417), .I1(n10601), .I2(n10580), .I3(port_id[3]), 
            .O(n11420));
    defparam n11417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10313 (.I0(port_id[2]), .I1(n8957), .I2(n8966), 
            .I3(port_id[3]), .O(n11411));
    defparam port_id_2__bdd_4_lut_10313.LUT_INIT = 16'he4aa;
    SB_LUT4 n11411_bdd_4_lut (.I0(n11411), .I1(n8933), .I2(n8921), .I3(port_id[3]), 
            .O(n11414));
    defparam n11411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10318 (.I0(port_id[0]), .I1(ram_s_58_2), 
            .I2(ram_s_59_2), .I3(port_id[1]), .O(n11405));
    defparam port_id_0__bdd_4_lut_10318.LUT_INIT = 16'he4aa;
    SB_LUT4 n11405_bdd_4_lut (.I0(n11405), .I1(ram_s_57_2), .I2(ram_s_56_2), 
            .I3(port_id[1]), .O(n11408));
    defparam n11405_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10308 (.I0(port_id[2]), .I1(n10319), .I2(n10352), 
            .I3(port_id[3]), .O(n11399));
    defparam port_id_2__bdd_4_lut_10308.LUT_INIT = 16'he4aa;
    SB_LUT4 n11399_bdd_4_lut (.I0(n11399), .I1(n10283), .I2(n10247), .I3(port_id[3]), 
            .O(n11402));
    defparam n11399_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10303 (.I0(port_id[0]), .I1(ram_s_174_5), 
            .I2(ram_s_175_5), .I3(port_id[1]), .O(n11393));
    defparam port_id_0__bdd_4_lut_10303.LUT_INIT = 16'he4aa;
    SB_LUT4 n11393_bdd_4_lut (.I0(n11393), .I1(ram_s_173_5), .I2(ram_s_172_5), 
            .I3(port_id[1]), .O(n11396));
    defparam n11393_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10293 (.I0(port_id[0]), .I1(ram_s_222_5), 
            .I2(ram_s_223_5), .I3(port_id[1]), .O(n11387));
    defparam port_id_0__bdd_4_lut_10293.LUT_INIT = 16'he4aa;
    SB_LUT4 n11387_bdd_4_lut (.I0(n11387), .I1(ram_s_221_5), .I2(ram_s_220_5), 
            .I3(port_id[1]), .O(n11390));
    defparam n11387_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10288 (.I0(port_id[0]), .I1(ram_s_98_5), 
            .I2(ram_s_99_5), .I3(port_id[1]), .O(n11381));
    defparam port_id_0__bdd_4_lut_10288.LUT_INIT = 16'he4aa;
    SB_LUT4 n11381_bdd_4_lut (.I0(n11381), .I1(ram_s_97_5), .I2(ram_s_96_5), 
            .I3(port_id[1]), .O(n11384));
    defparam n11381_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1519_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_109_7), .O(n1767));   // src/ram.vhd(68[19:45])
    defparam i1519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1518_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_109_6), .O(n1766));   // src/ram.vhd(68[19:45])
    defparam i1518_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_2__bdd_4_lut_10298 (.I0(port_id[2]), .I1(n9467), .I2(n9752), 
            .I3(port_id[3]), .O(n11375));
    defparam port_id_2__bdd_4_lut_10298.LUT_INIT = 16'he4aa;
    SB_LUT4 n11375_bdd_4_lut (.I0(n11375), .I1(n11366), .I2(n11330), .I3(port_id[3]), 
            .O(n10562));
    defparam n11375_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10283 (.I0(port_id[0]), .I1(ram_s_62_2), 
            .I2(ram_s_63_2), .I3(port_id[1]), .O(n11369));
    defparam port_id_0__bdd_4_lut_10283.LUT_INIT = 16'he4aa;
    SB_LUT4 n11369_bdd_4_lut (.I0(n11369), .I1(ram_s_61_2), .I2(ram_s_60_2), 
            .I3(port_id[1]), .O(n11372));
    defparam n11369_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10273 (.I0(port_id[0]), .I1(ram_s_22_5), 
            .I2(ram_s_23_5), .I3(port_id[1]), .O(n11363));
    defparam port_id_0__bdd_4_lut_10273.LUT_INIT = 16'he4aa;
    SB_LUT4 n11363_bdd_4_lut (.I0(n11363), .I1(ram_s_21_5), .I2(ram_s_20_5), 
            .I3(port_id[1]), .O(n11366));
    defparam n11363_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_10338 (.I0(port_id[1]), .I1(n9639), .I2(n9640), 
            .I3(port_id[2]), .O(n11357));
    defparam port_id_1__bdd_4_lut_10338.LUT_INIT = 16'he4aa;
    SB_LUT4 n11357_bdd_4_lut (.I0(n11357), .I1(n9622), .I2(n9621), .I3(port_id[2]), 
            .O(n11360));
    defparam n11357_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10268 (.I0(port_id[0]), .I1(ram_s_50_3), 
            .I2(ram_s_51_3), .I3(port_id[1]), .O(n11351));
    defparam port_id_0__bdd_4_lut_10268.LUT_INIT = 16'he4aa;
    SB_LUT4 n11351_bdd_4_lut (.I0(n11351), .I1(ram_s_49_3), .I2(ram_s_48_3), 
            .I3(port_id[1]), .O(n11354));
    defparam n11351_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_10263 (.I0(port_id[1]), .I1(n9441), .I2(n9442), 
            .I3(port_id[2]), .O(n11333));
    defparam port_id_1__bdd_4_lut_10263.LUT_INIT = 16'he4aa;
    SB_LUT4 n11333_bdd_4_lut (.I0(n11333), .I1(n9424), .I2(n9423), .I3(port_id[2]), 
            .O(n11336));
    defparam n11333_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2032_3_lut_4_lut (.I0(n228), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_174_0), .O(n2280));   // src/ram.vhd(68[19:45])
    defparam i2032_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10258 (.I0(port_id[0]), .I1(ram_s_18_5), 
            .I2(ram_s_19_5), .I3(port_id[1]), .O(n11327));
    defparam port_id_0__bdd_4_lut_10258.LUT_INIT = 16'he4aa;
    SB_LUT4 n11327_bdd_4_lut (.I0(n11327), .I1(ram_s_17_5), .I2(ram_s_16_5), 
            .I3(port_id[1]), .O(n11330));
    defparam n11327_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_10243 (.I0(port_id[1]), .I1(n10068), .I2(n10069), 
            .I3(port_id[2]), .O(n11321));
    defparam port_id_1__bdd_4_lut_10243.LUT_INIT = 16'he4aa;
    SB_LUT4 n11321_bdd_4_lut (.I0(n11321), .I1(n10060), .I2(n10059), .I3(port_id[2]), 
            .O(n11324));
    defparam n11321_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1517_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_109_5), .O(n1765));   // src/ram.vhd(68[19:45])
    defparam i1517_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10238 (.I0(port_id[0]), .I1(ram_s_66_2), 
            .I2(ram_s_67_2), .I3(port_id[1]), .O(n11309));
    defparam port_id_0__bdd_4_lut_10238.LUT_INIT = 16'he4aa;
    SB_LUT4 n11309_bdd_4_lut (.I0(n11309), .I1(ram_s_65_2), .I2(ram_s_64_2), 
            .I3(port_id[1]), .O(n11312));
    defparam n11309_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10224 (.I0(port_id[0]), .I1(ram_s_154_3), 
            .I2(ram_s_155_3), .I3(port_id[1]), .O(n11297));
    defparam port_id_0__bdd_4_lut_10224.LUT_INIT = 16'he4aa;
    SB_LUT4 n11297_bdd_4_lut (.I0(n11297), .I1(ram_s_153_3), .I2(ram_s_152_3), 
            .I3(port_id[1]), .O(n9794));
    defparam n11297_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1516_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_109_4), .O(n1764));   // src/ram.vhd(68[19:45])
    defparam i1516_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10214 (.I0(port_id[0]), .I1(ram_s_46_1), 
            .I2(ram_s_47_1), .I3(port_id[1]), .O(n11291));
    defparam port_id_0__bdd_4_lut_10214.LUT_INIT = 16'he4aa;
    SB_LUT4 n11291_bdd_4_lut (.I0(n11291), .I1(ram_s_45_1), .I2(ram_s_44_1), 
            .I3(port_id[1]), .O(n11294));
    defparam n11291_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10209 (.I0(port_id[0]), .I1(ram_s_46_0), 
            .I2(ram_s_47_0), .I3(port_id[1]), .O(n11285));
    defparam port_id_0__bdd_4_lut_10209.LUT_INIT = 16'he4aa;
    SB_LUT4 n11285_bdd_4_lut (.I0(n11285), .I1(ram_s_45_0), .I2(ram_s_44_0), 
            .I3(port_id[1]), .O(n11288));
    defparam n11285_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i354_2_lut_3_lut (.I0(n97_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n212));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i354_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 port_id_0__bdd_4_lut_10204 (.I0(port_id[0]), .I1(ram_s_70_2), 
            .I2(ram_s_71_2), .I3(port_id[1]), .O(n11279));
    defparam port_id_0__bdd_4_lut_10204.LUT_INIT = 16'he4aa;
    SB_LUT4 n11279_bdd_4_lut (.I0(n11279), .I1(ram_s_69_2), .I2(ram_s_68_2), 
            .I3(port_id[1]), .O(n11282));
    defparam n11279_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10199 (.I0(port_id[0]), .I1(ram_s_50_1), 
            .I2(ram_s_51_1), .I3(port_id[1]), .O(n11267));
    defparam port_id_0__bdd_4_lut_10199.LUT_INIT = 16'he4aa;
    SB_LUT4 n11267_bdd_4_lut (.I0(n11267), .I1(ram_s_49_1), .I2(ram_s_48_1), 
            .I3(port_id[1]), .O(n11270));
    defparam n11267_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1515_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_109_3), .O(n1763));   // src/ram.vhd(68[19:45])
    defparam i1515_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_1__bdd_4_lut_10233 (.I0(port_id[1]), .I1(n9234), .I2(n9235), 
            .I3(port_id[2]), .O(n11255));
    defparam port_id_1__bdd_4_lut_10233.LUT_INIT = 16'he4aa;
    SB_LUT4 n11255_bdd_4_lut (.I0(n11255), .I1(n9217), .I2(n9216), .I3(port_id[2]), 
            .O(n11258));
    defparam n11255_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10190 (.I0(port_id[0]), .I1(ram_s_222_7), 
            .I2(ram_s_223_7), .I3(port_id[1]), .O(n11249));
    defparam port_id_0__bdd_4_lut_10190.LUT_INIT = 16'he4aa;
    SB_LUT4 n11249_bdd_4_lut (.I0(n11249), .I1(ram_s_221_7), .I2(ram_s_220_7), 
            .I3(port_id[1]), .O(n11252));
    defparam n11249_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10278 (.I0(port_id[2]), .I1(n9110), .I2(n9122), 
            .I3(port_id[3]), .O(n11243));
    defparam port_id_2__bdd_4_lut_10278.LUT_INIT = 16'he4aa;
    SB_LUT4 n11243_bdd_4_lut (.I0(n11243), .I1(n9107), .I2(n9098), .I3(port_id[3]), 
            .O(n11246));
    defparam n11243_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_10402 (.I0(port_id[4]), .I1(n10592), .I2(n10628), 
            .I3(port_id[5]), .O(n11237));
    defparam port_id_4__bdd_4_lut_10402.LUT_INIT = 16'he4aa;
    SB_LUT4 n11237_bdd_4_lut (.I0(n11237), .I1(n10562), .I2(n10529), .I3(port_id[5]), 
            .O(n11240));
    defparam n11237_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i353_2_lut_3_lut (.I0(n97_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n84));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i353_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1514_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_109_2), .O(n1762));   // src/ram.vhd(68[19:45])
    defparam i1514_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i352_2_lut_3_lut (.I0(n95_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n213));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i352_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i351_2_lut_3_lut (.I0(n95_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n85));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i351_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i350_2_lut_3_lut (.I0(n93_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n214));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i350_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i349_2_lut_3_lut (.I0(n93_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n86));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i349_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2007_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_170_7), .O(n2255));   // src/ram.vhd(68[19:45])
    defparam i2007_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1513_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_109_1), .O(n1761));   // src/ram.vhd(68[19:45])
    defparam i1513_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1512_3_lut_4_lut (.I0(n225_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_109_0), .O(n1760));   // src/ram.vhd(68[19:45])
    defparam i1512_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2487_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_230_7), .O(n2735));   // src/ram.vhd(68[19:45])
    defparam i2487_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2006_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_170_6), .O(n2254));   // src/ram.vhd(68[19:45])
    defparam i2006_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2005_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_170_5), .O(n2253));   // src/ram.vhd(68[19:45])
    defparam i2005_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2004_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_170_4), .O(n2252));   // src/ram.vhd(68[19:45])
    defparam i2004_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2486_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_230_6), .O(n2734));   // src/ram.vhd(68[19:45])
    defparam i2486_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2485_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_230_5), .O(n2733));   // src/ram.vhd(68[19:45])
    defparam i2485_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2003_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_170_3), .O(n2251));   // src/ram.vhd(68[19:45])
    defparam i2003_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2484_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_230_4), .O(n2732));   // src/ram.vhd(68[19:45])
    defparam i2484_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2002_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_170_2), .O(n2250));   // src/ram.vhd(68[19:45])
    defparam i2002_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2483_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_230_3), .O(n2731));   // src/ram.vhd(68[19:45])
    defparam i2483_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2001_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_170_1), .O(n2249));   // src/ram.vhd(68[19:45])
    defparam i2001_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2482_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_230_2), .O(n2730));   // src/ram.vhd(68[19:45])
    defparam i2482_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2481_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_230_1), .O(n2729));   // src/ram.vhd(68[19:45])
    defparam i2481_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i199_2_lut (.I0(n71_adj_842), .I1(port_id[6]), 
            .I2(wea[0]), .I3(wea[0]), .O(n199_adj_843));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2480_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_230_0), .O(n2728));   // src/ram.vhd(68[19:45])
    defparam i2480_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2000_3_lut_4_lut (.I0(n220_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_170_0), .O(n2248));   // src/ram.vhd(68[19:45])
    defparam i2000_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1999_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_169_7), .O(n2247));   // src/ram.vhd(68[19:45])
    defparam i1999_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1998_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_169_6), .O(n2246));   // src/ram.vhd(68[19:45])
    defparam i1998_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1997_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_169_5), .O(n2245));   // src/ram.vhd(68[19:45])
    defparam i1997_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1996_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_169_4), .O(n2244));   // src/ram.vhd(68[19:45])
    defparam i1996_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1995_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_169_3), .O(n2243));   // src/ram.vhd(68[19:45])
    defparam i1995_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1994_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_169_2), .O(n2242));   // src/ram.vhd(68[19:45])
    defparam i1994_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1993_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_169_1), .O(n2241));   // src/ram.vhd(68[19:45])
    defparam i1993_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_2__bdd_4_lut_11129 (.I0(port_id[2]), .I1(n9629), .I2(n9701), 
            .I3(port_id[3]), .O(n12311));
    defparam port_id_2__bdd_4_lut_11129.LUT_INIT = 16'he4aa;
    SB_LUT4 n12311_bdd_4_lut (.I0(n12311), .I1(n9557), .I2(n9491), .I3(port_id[3]), 
            .O(n12314));
    defparam n12311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10436 (.I0(port_id[2]), .I1(n9650), .I2(n9680), 
            .I3(port_id[3]), .O(n11555));
    defparam port_id_2__bdd_4_lut_10436.LUT_INIT = 16'he4aa;
    SB_LUT4 n11555_bdd_4_lut (.I0(n11555), .I1(n9605), .I2(n9584), .I3(port_id[3]), 
            .O(n11558));
    defparam n11555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10870 (.I0(port_id[0]), .I1(ram_s_174_1), 
            .I2(ram_s_175_1), .I3(port_id[1]), .O(n12083));
    defparam port_id_0__bdd_4_lut_10870.LUT_INIT = 16'he4aa;
    SB_LUT4 n12083_bdd_4_lut (.I0(n12083), .I1(ram_s_173_1), .I2(ram_s_172_1), 
            .I3(port_id[1]), .O(n12086));
    defparam n12083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11060 (.I0(port_id[0]), .I1(ram_s_174_6), 
            .I2(ram_s_175_6), .I3(port_id[1]), .O(n12305));
    defparam port_id_0__bdd_4_lut_11060.LUT_INIT = 16'he4aa;
    SB_LUT4 n12305_bdd_4_lut (.I0(n12305), .I1(ram_s_173_6), .I2(ram_s_172_6), 
            .I3(port_id[1]), .O(n12308));
    defparam n12305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1992_3_lut_4_lut (.I0(n218_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_169_0), .O(n2240));   // src/ram.vhd(68[19:45])
    defparam i1992_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1511_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_108_7), .O(n1759));   // src/ram.vhd(68[19:45])
    defparam i1511_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i201_2_lut (.I0(n73), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n201));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1510_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_108_6), .O(n1758));   // src/ram.vhd(68[19:45])
    defparam i1510_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1509_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_108_5), .O(n1757));   // src/ram.vhd(68[19:45])
    defparam i1509_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i203_2_lut (.I0(n75), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n203));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1508_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_108_4), .O(n1756));   // src/ram.vhd(68[19:45])
    defparam i1508_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i344_2_lut_3_lut (.I0(n87), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n217));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i344_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i343_2_lut_3_lut (.I0(n87), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n89));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i343_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i342_2_lut_3_lut (.I0(n85_adj_845), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n218));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i342_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i341_2_lut_3_lut (.I0(n85_adj_845), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n90));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i341_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1507_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_108_3), .O(n1755));   // src/ram.vhd(68[19:45])
    defparam i1507_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i205_2_lut (.I0(n77), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n205));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1506_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_108_2), .O(n1754));   // src/ram.vhd(68[19:45])
    defparam i1506_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i340_2_lut_3_lut (.I0(n83), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n219));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i340_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i339_2_lut_3_lut (.I0(n83), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n91));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i339_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i338_2_lut_3_lut (.I0(n81), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n220));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i338_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i337_2_lut_3_lut (.I0(n81), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n92));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i337_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i336_2_lut_3_lut (.I0(n79), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n221));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i336_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1505_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_108_1), .O(n1753));   // src/ram.vhd(68[19:45])
    defparam i1505_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1504_3_lut_4_lut (.I0(n223_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_108_0), .O(n1752));   // src/ram.vhd(68[19:45])
    defparam i1504_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i207_2_lut (.I0(n79), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n207));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 EnabledDecoder_2_i335_2_lut_3_lut (.I0(n79), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n93));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i335_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i334_2_lut_3_lut (.I0(n77), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n222));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i334_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i2479_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_229_7), .O(n2727));   // src/ram.vhd(68[19:45])
    defparam i2479_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i209_2_lut (.I0(n81), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n209));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 EnabledDecoder_2_i333_2_lut_3_lut (.I0(n77), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n94));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i333_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2478_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_229_6), .O(n2726));   // src/ram.vhd(68[19:45])
    defparam i2478_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2477_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_229_5), .O(n2725));   // src/ram.vhd(68[19:45])
    defparam i2477_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i332_2_lut_3_lut (.I0(n75), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n223));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i332_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i2476_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_229_4), .O(n2724));   // src/ram.vhd(68[19:45])
    defparam i2476_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i331_2_lut_3_lut (.I0(n75), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n95));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i331_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i330_2_lut_3_lut (.I0(n73), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n224));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i330_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i2321_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_210_1), .O(n2569));   // src/ram.vhd(68[19:45])
    defparam i2321_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i211_2_lut (.I0(n83), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n211));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 EnabledDecoder_2_i329_2_lut_3_lut (.I0(n73), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n96));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i329_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2475_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_229_3), .O(n2723));   // src/ram.vhd(68[19:45])
    defparam i2475_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2474_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_229_2), .O(n2722));   // src/ram.vhd(68[19:45])
    defparam i2474_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i328_2_lut_3_lut (.I0(n71_adj_842), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n225));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i328_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i213_2_lut (.I0(n85_adj_845), .I1(port_id[6]), 
            .I2(wea[0]), .I3(wea[0]), .O(n213_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 EnabledDecoder_2_i327_2_lut_3_lut (.I0(n71_adj_842), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n97));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i327_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2473_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_229_1), .O(n2721));   // src/ram.vhd(68[19:45])
    defparam i2473_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1919_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_159_7), .O(n2167));   // src/ram.vhd(68[19:45])
    defparam i1919_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1918_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_159_6), .O(n2166));   // src/ram.vhd(68[19:45])
    defparam i1918_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1917_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_159_5), .O(n2165));   // src/ram.vhd(68[19:45])
    defparam i1917_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2472_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_229_0), .O(n2720));   // src/ram.vhd(68[19:45])
    defparam i2472_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i215_2_lut (.I0(n87), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n215));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1916_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_159_4), .O(n2164));   // src/ram.vhd(68[19:45])
    defparam i1916_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1915_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_159_3), .O(n2163));   // src/ram.vhd(68[19:45])
    defparam i1915_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1914_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_159_2), .O(n2162));   // src/ram.vhd(68[19:45])
    defparam i1914_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1913_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_159_1), .O(n2161));   // src/ram.vhd(68[19:45])
    defparam i1913_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1912_3_lut_4_lut (.I0(n198), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_159_0), .O(n2160));   // src/ram.vhd(68[19:45])
    defparam i1912_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1911_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_158_7), .O(n2159));   // src/ram.vhd(68[19:45])
    defparam i1911_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1910_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_158_6), .O(n2158));   // src/ram.vhd(68[19:45])
    defparam i1910_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1909_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_158_5), .O(n2157));   // src/ram.vhd(68[19:45])
    defparam i1909_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2471_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_228_7), .O(n2719));   // src/ram.vhd(68[19:45])
    defparam i2471_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1908_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_158_4), .O(n2156));   // src/ram.vhd(68[19:45])
    defparam i1908_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2470_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_228_6), .O(n2718));   // src/ram.vhd(68[19:45])
    defparam i2470_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1907_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_158_3), .O(n2155));   // src/ram.vhd(68[19:45])
    defparam i1907_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1906_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_158_2), .O(n2154));   // src/ram.vhd(68[19:45])
    defparam i1906_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2469_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_228_5), .O(n2717));   // src/ram.vhd(68[19:45])
    defparam i2469_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i221_2_lut (.I0(n93_c), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n221_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1905_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_158_1), .O(n2153));   // src/ram.vhd(68[19:45])
    defparam i1905_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1904_3_lut_4_lut (.I0(n196), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_158_0), .O(n2152));   // src/ram.vhd(68[19:45])
    defparam i1904_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i650_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_10_2), .O(n898));   // src/ram.vhd(68[19:45])
    defparam i650_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i647_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_10_3), .O(n895));   // src/ram.vhd(68[19:45])
    defparam i647_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i446_447 (.Q(ram_s_18_0), .C(CLK_3P3_MHZ_c), .D(n921));   // src/ram.vhd(56[12:17])
    SB_DFF i443_444 (.Q(ram_s_17_7), .C(CLK_3P3_MHZ_c), .D(n920));   // src/ram.vhd(56[12:17])
    SB_DFF i449_450 (.Q(ram_s_18_1), .C(CLK_3P3_MHZ_c), .D(n919));   // src/ram.vhd(56[12:17])
    SB_DFF i347_348 (.Q(ram_s_13_7), .C(CLK_3P3_MHZ_c), .D(n918));   // src/ram.vhd(56[12:17])
    SB_DFF i350_351 (.Q(ram_s_14_0), .C(CLK_3P3_MHZ_c), .D(n917));   // src/ram.vhd(56[12:17])
    SB_DFF i353_354 (.Q(ram_s_14_1), .C(CLK_3P3_MHZ_c), .D(n916));   // src/ram.vhd(56[12:17])
    SB_DFF i518_519 (.Q(ram_s_21_0), .C(CLK_3P3_MHZ_c), .D(n915));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2468_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_228_4), .O(n2716));   // src/ram.vhd(68[19:45])
    defparam i2468_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i648_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_10_0), .O(n896));   // src/ram.vhd(68[19:45])
    defparam i648_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2467_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_228_3), .O(n2715));   // src/ram.vhd(68[19:45])
    defparam i2467_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i223_2_lut (.I0(n95_c), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n223_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i646_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_10_1), .O(n894));   // src/ram.vhd(68[19:45])
    defparam i646_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2466_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_228_2), .O(n2714));   // src/ram.vhd(68[19:45])
    defparam i2466_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i662_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_10_7), .O(n910));   // src/ram.vhd(68[19:45])
    defparam i662_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i700_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_10_6), .O(n948));   // src/ram.vhd(68[19:45])
    defparam i700_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2465_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_228_1), .O(n2713));   // src/ram.vhd(68[19:45])
    defparam i2465_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i225_2_lut (.I0(n97_c), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n225_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2464_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_228_0), .O(n2712));   // src/ram.vhd(68[19:45])
    defparam i2464_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i701_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_10_5), .O(n949));   // src/ram.vhd(68[19:45])
    defparam i701_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i638_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_10_4), .O(n886));   // src/ram.vhd(68[19:45])
    defparam i638_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2320_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_210_0), .O(n2568));   // src/ram.vhd(68[19:45])
    defparam i2320_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10123 (.I0(port_id[0]), .I1(ram_s_50_2), 
            .I2(ram_s_51_2), .I3(port_id[1]), .O(n11177));
    defparam port_id_0__bdd_4_lut_10123.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i219_2_lut_3_lut_4_lut (.I0(n27), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n219_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i219_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 n11177_bdd_4_lut (.I0(n11177), .I1(ram_s_49_2), .I2(ram_s_48_2), 
            .I3(port_id[1]), .O(n11180));
    defparam n11177_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i220_2_lut_3_lut_4_lut (.I0(n27), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n220_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i220_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1503_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_107_7), .O(n1751));   // src/ram.vhd(68[19:45])
    defparam i1503_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1311_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_83_7), .O(n1559));   // src/ram.vhd(68[19:45])
    defparam i1311_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1502_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_107_6), .O(n1750));   // src/ram.vhd(68[19:45])
    defparam i1502_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i11_2_lut_3_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[1]), .I3(wea[0]), .O(n11));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i11_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i15_2_lut_3_lut_4_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[2]), .I3(port_id[1]), .O(n15));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i15_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1501_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_107_5), .O(n1749));   // src/ram.vhd(68[19:45])
    defparam i1501_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1500_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_107_4), .O(n1748));   // src/ram.vhd(68[19:45])
    defparam i1500_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i229_2_lut (.I0(n101), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n229));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 EnabledDecoder_2_i16_2_lut_3_lut_4_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[2]), .I3(port_id[1]), .O(n16));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i16_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1499_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_107_3), .O(n1747));   // src/ram.vhd(68[19:45])
    defparam i1499_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1498_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_107_2), .O(n1746));   // src/ram.vhd(68[19:45])
    defparam i1498_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1497_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_107_1), .O(n1745));   // src/ram.vhd(68[19:45])
    defparam i1497_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1496_3_lut_4_lut (.I0(n221_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_107_0), .O(n1744));   // src/ram.vhd(68[19:45])
    defparam i1496_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2463_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_227_7), .O(n2711));   // src/ram.vhd(68[19:45])
    defparam i2463_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2462_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_227_6), .O(n2710));   // src/ram.vhd(68[19:45])
    defparam i2462_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1310_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_83_6), .O(n1558));   // src/ram.vhd(68[19:45])
    defparam i1310_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2461_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_227_5), .O(n2709));   // src/ram.vhd(68[19:45])
    defparam i2461_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1309_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_83_5), .O(n1557));   // src/ram.vhd(68[19:45])
    defparam i1309_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2460_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_227_4), .O(n2708));   // src/ram.vhd(68[19:45])
    defparam i2460_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1308_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_83_4), .O(n1556));   // src/ram.vhd(68[19:45])
    defparam i1308_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2459_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_227_3), .O(n2707));   // src/ram.vhd(68[19:45])
    defparam i2459_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2458_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_227_2), .O(n2706));   // src/ram.vhd(68[19:45])
    defparam i2458_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2457_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_227_1), .O(n2705));   // src/ram.vhd(68[19:45])
    defparam i2457_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1307_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_83_3), .O(n1555));   // src/ram.vhd(68[19:45])
    defparam i1307_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2456_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_227_0), .O(n2704));   // src/ram.vhd(68[19:45])
    defparam i2456_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1495_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_106_7), .O(n1743));   // src/ram.vhd(68[19:45])
    defparam i1495_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i249_2_lut (.I0(n121_c), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n249_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1494_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_106_6), .O(n1742));   // src/ram.vhd(68[19:45])
    defparam i1494_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1903_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_157_7), .O(n2151));   // src/ram.vhd(68[19:45])
    defparam i1903_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1902_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_157_6), .O(n2150));   // src/ram.vhd(68[19:45])
    defparam i1902_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1493_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_106_5), .O(n1741));   // src/ram.vhd(68[19:45])
    defparam i1493_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1901_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_157_5), .O(n2149));   // src/ram.vhd(68[19:45])
    defparam i1901_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1492_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_106_4), .O(n1740));   // src/ram.vhd(68[19:45])
    defparam i1492_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1491_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_106_3), .O(n1739));   // src/ram.vhd(68[19:45])
    defparam i1491_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1490_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_106_2), .O(n1738));   // src/ram.vhd(68[19:45])
    defparam i1490_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i251_2_lut (.I0(n123_c), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n251_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1900_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_157_4), .O(n2148));   // src/ram.vhd(68[19:45])
    defparam i1900_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1489_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_106_1), .O(n1737));   // src/ram.vhd(68[19:45])
    defparam i1489_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1899_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_157_3), .O(n2147));   // src/ram.vhd(68[19:45])
    defparam i1899_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1488_3_lut_4_lut (.I0(n219_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_106_0), .O(n1736));   // src/ram.vhd(68[19:45])
    defparam i1488_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2455_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_226_7), .O(n2703));   // src/ram.vhd(68[19:45])
    defparam i2455_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1898_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_157_2), .O(n2146));   // src/ram.vhd(68[19:45])
    defparam i1898_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2454_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_226_6), .O(n2702));   // src/ram.vhd(68[19:45])
    defparam i2454_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2453_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_226_5), .O(n2701));   // src/ram.vhd(68[19:45])
    defparam i2453_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1897_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_157_1), .O(n2145));   // src/ram.vhd(68[19:45])
    defparam i1897_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2452_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_226_4), .O(n2700));   // src/ram.vhd(68[19:45])
    defparam i2452_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2451_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_226_3), .O(n2699));   // src/ram.vhd(68[19:45])
    defparam i2451_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1896_3_lut_4_lut (.I0(n194_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_157_0), .O(n2144));   // src/ram.vhd(68[19:45])
    defparam i1896_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2450_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_226_2), .O(n2698));   // src/ram.vhd(68[19:45])
    defparam i2450_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2449_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_226_1), .O(n2697));   // src/ram.vhd(68[19:45])
    defparam i2449_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2448_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_226_0), .O(n2696));   // src/ram.vhd(68[19:45])
    defparam i2448_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i259_2_lut (.I0(n131), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n259));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1895_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_156_7), .O(n2143));   // src/ram.vhd(68[19:45])
    defparam i1895_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1894_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_156_6), .O(n2142));   // src/ram.vhd(68[19:45])
    defparam i1894_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i37_2_lut (.I0(n21), .I1(port_id[3]), .I2(wea[0]), 
            .I3(wea[0]), .O(n37));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i37_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1893_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_156_5), .O(n2141));   // src/ram.vhd(68[19:45])
    defparam i1893_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1487_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_105_7), .O(n1735));   // src/ram.vhd(68[19:45])
    defparam i1487_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1486_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_105_6), .O(n1734));   // src/ram.vhd(68[19:45])
    defparam i1486_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1892_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_156_4), .O(n2140));   // src/ram.vhd(68[19:45])
    defparam i1892_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1891_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_156_3), .O(n2139));   // src/ram.vhd(68[19:45])
    defparam i1891_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1306_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_83_2), .O(n1554));   // src/ram.vhd(68[19:45])
    defparam i1306_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1485_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_105_5), .O(n1733));   // src/ram.vhd(68[19:45])
    defparam i1485_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i261_2_lut (.I0(n133), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n261));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1890_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_156_2), .O(n2138));   // src/ram.vhd(68[19:45])
    defparam i1890_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1889_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_156_1), .O(n2137));   // src/ram.vhd(68[19:45])
    defparam i1889_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1484_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_105_4), .O(n1732));   // src/ram.vhd(68[19:45])
    defparam i1484_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1305_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_83_1), .O(n1553));   // src/ram.vhd(68[19:45])
    defparam i1305_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1888_3_lut_4_lut (.I0(n192_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_156_0), .O(n2136));   // src/ram.vhd(68[19:45])
    defparam i1888_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1483_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_105_3), .O(n1731));   // src/ram.vhd(68[19:45])
    defparam i1483_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2301_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_207_5), .O(n2549));   // src/ram.vhd(68[19:45])
    defparam i2301_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1482_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_105_2), .O(n1730));   // src/ram.vhd(68[19:45])
    defparam i1482_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1481_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_105_1), .O(n1729));   // src/ram.vhd(68[19:45])
    defparam i1481_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1480_3_lut_4_lut (.I0(n217_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_105_0), .O(n1728));   // src/ram.vhd(68[19:45])
    defparam i1480_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2300_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_207_4), .O(n2548));   // src/ram.vhd(68[19:45])
    defparam i2300_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2447_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_225_7), .O(n2695));   // src/ram.vhd(68[19:45])
    defparam i2447_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1887_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_155_7), .O(n2135));   // src/ram.vhd(68[19:45])
    defparam i1887_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1886_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_155_6), .O(n2134));   // src/ram.vhd(68[19:45])
    defparam i1886_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1885_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_155_5), .O(n2133));   // src/ram.vhd(68[19:45])
    defparam i1885_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1304_3_lut_4_lut (.I0(n173), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_83_0), .O(n1552));   // src/ram.vhd(68[19:45])
    defparam i1304_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_4__bdd_4_lut_10165 (.I0(port_id[4]), .I1(n10250), .I2(n8813), 
            .I3(port_id[5]), .O(n11171));
    defparam port_id_4__bdd_4_lut_10165.LUT_INIT = 16'he4aa;
    SB_LUT4 i2446_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_225_6), .O(n2694));   // src/ram.vhd(68[19:45])
    defparam i2446_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1884_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_155_4), .O(n2132));   // src/ram.vhd(68[19:45])
    defparam i1884_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1883_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_155_3), .O(n2131));   // src/ram.vhd(68[19:45])
    defparam i1883_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1882_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_155_2), .O(n2130));   // src/ram.vhd(68[19:45])
    defparam i1882_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2445_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_225_5), .O(n2693));   // src/ram.vhd(68[19:45])
    defparam i2445_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2444_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_225_4), .O(n2692));   // src/ram.vhd(68[19:45])
    defparam i2444_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1881_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_155_1), .O(n2129));   // src/ram.vhd(68[19:45])
    defparam i1881_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1880_3_lut_4_lut (.I0(n190_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_155_0), .O(n2128));   // src/ram.vhd(68[19:45])
    defparam i1880_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2443_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_225_3), .O(n2691));   // src/ram.vhd(68[19:45])
    defparam i2443_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i172_2_lut_3_lut (.I0(n43), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n172));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i172_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 n11171_bdd_4_lut (.I0(n11171), .I1(n8798), .I2(n8855), .I3(port_id[5]), 
            .O(n11174));
    defparam n11171_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2442_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_225_2), .O(n2690));   // src/ram.vhd(68[19:45])
    defparam i2442_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i171_2_lut_3_lut (.I0(n43), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n171));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i171_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2441_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_225_1), .O(n2689));   // src/ram.vhd(68[19:45])
    defparam i2441_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2440_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_225_0), .O(n2688));   // src/ram.vhd(68[19:45])
    defparam i2440_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1303_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_82_7), .O(n1551));   // src/ram.vhd(68[19:45])
    defparam i1303_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1302_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_82_6), .O(n1550));   // src/ram.vhd(68[19:45])
    defparam i1302_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2299_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_207_3), .O(n2547));   // src/ram.vhd(68[19:45])
    defparam i2299_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1479_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_104_7), .O(n1727));   // src/ram.vhd(68[19:45])
    defparam i1479_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1478_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_104_6), .O(n1726));   // src/ram.vhd(68[19:45])
    defparam i1478_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1477_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_104_5), .O(n1725));   // src/ram.vhd(68[19:45])
    defparam i1477_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1476_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_104_4), .O(n1724));   // src/ram.vhd(68[19:45])
    defparam i1476_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1475_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_104_3), .O(n1723));   // src/ram.vhd(68[19:45])
    defparam i1475_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1474_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_104_2), .O(n1722));   // src/ram.vhd(68[19:45])
    defparam i1474_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1473_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_104_1), .O(n1721));   // src/ram.vhd(68[19:45])
    defparam i1473_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1472_3_lut_4_lut (.I0(n215), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_104_0), .O(n1720));   // src/ram.vhd(68[19:45])
    defparam i1472_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2439_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_224_7), .O(n2687));   // src/ram.vhd(68[19:45])
    defparam i2439_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2438_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_224_6), .O(n2686));   // src/ram.vhd(68[19:45])
    defparam i2438_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2437_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_224_5), .O(n2685));   // src/ram.vhd(68[19:45])
    defparam i2437_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2436_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_224_4), .O(n2684));   // src/ram.vhd(68[19:45])
    defparam i2436_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1879_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_154_7), .O(n2127));   // src/ram.vhd(68[19:45])
    defparam i1879_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2298_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_207_2), .O(n2546));   // src/ram.vhd(68[19:45])
    defparam i2298_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2435_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_224_3), .O(n2683));   // src/ram.vhd(68[19:45])
    defparam i2435_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1301_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_82_5), .O(n1549));   // src/ram.vhd(68[19:45])
    defparam i1301_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2434_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_224_2), .O(n2682));   // src/ram.vhd(68[19:45])
    defparam i2434_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2433_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_224_1), .O(n2681));   // src/ram.vhd(68[19:45])
    defparam i2433_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1878_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_154_6), .O(n2126));   // src/ram.vhd(68[19:45])
    defparam i1878_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1877_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_154_5), .O(n2125));   // src/ram.vhd(68[19:45])
    defparam i1877_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2432_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_224_0), .O(n2680));   // src/ram.vhd(68[19:45])
    defparam i2432_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1876_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_154_4), .O(n2124));   // src/ram.vhd(68[19:45])
    defparam i1876_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1875_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_154_3), .O(n2123));   // src/ram.vhd(68[19:45])
    defparam i1875_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1471_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_103_7), .O(n1719));   // src/ram.vhd(68[19:45])
    defparam i1471_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1874_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_154_2), .O(n2122));   // src/ram.vhd(68[19:45])
    defparam i1874_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1873_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_154_1), .O(n2121));   // src/ram.vhd(68[19:45])
    defparam i1873_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1872_3_lut_4_lut (.I0(n188_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_154_0), .O(n2120));   // src/ram.vhd(68[19:45])
    defparam i1872_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1470_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_103_6), .O(n1718));   // src/ram.vhd(68[19:45])
    defparam i1470_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1871_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_153_7), .O(n2119));   // src/ram.vhd(68[19:45])
    defparam i1871_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1469_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_103_5), .O(n1717));   // src/ram.vhd(68[19:45])
    defparam i1469_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1870_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_153_6), .O(n2118));   // src/ram.vhd(68[19:45])
    defparam i1870_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1468_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_103_4), .O(n1716));   // src/ram.vhd(68[19:45])
    defparam i1468_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1467_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_103_3), .O(n1715));   // src/ram.vhd(68[19:45])
    defparam i1467_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1869_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_153_5), .O(n2117));   // src/ram.vhd(68[19:45])
    defparam i1869_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1868_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_153_4), .O(n2116));   // src/ram.vhd(68[19:45])
    defparam i1868_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1466_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_103_2), .O(n1714));   // src/ram.vhd(68[19:45])
    defparam i1466_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1867_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_153_3), .O(n2115));   // src/ram.vhd(68[19:45])
    defparam i1867_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1866_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_153_2), .O(n2114));   // src/ram.vhd(68[19:45])
    defparam i1866_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1465_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_103_1), .O(n1713));   // src/ram.vhd(68[19:45])
    defparam i1465_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1865_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_153_1), .O(n2113));   // src/ram.vhd(68[19:45])
    defparam i1865_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1864_3_lut_4_lut (.I0(n186_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_153_0), .O(n2112));   // src/ram.vhd(68[19:45])
    defparam i1864_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1464_3_lut_4_lut (.I0(n213_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_103_0), .O(n1712));   // src/ram.vhd(68[19:45])
    defparam i1464_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2431_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_223_7), .O(n2679));   // src/ram.vhd(68[19:45])
    defparam i2431_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2430_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_223_6), .O(n2678));   // src/ram.vhd(68[19:45])
    defparam i2430_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8462_3_lut (.I0(n13172), .I1(n14480), .I2(port_id[7]), .I3(wea[0]), 
            .O(spm_ram_data[0]));
    defparam i8462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7925_3_lut (.I0(n11810), .I1(n14198), .I2(port_id[7]), .I3(wea[0]), 
            .O(spm_ram_data[7]));
    defparam i7925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2429_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_223_5), .O(n2677));   // src/ram.vhd(68[19:45])
    defparam i2429_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2428_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_223_4), .O(n2676));   // src/ram.vhd(68[19:45])
    defparam i2428_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2427_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_223_3), .O(n2675));   // src/ram.vhd(68[19:45])
    defparam i2427_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2426_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_223_2), .O(n2674));   // src/ram.vhd(68[19:45])
    defparam i2426_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2425_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_223_1), .O(n2673));   // src/ram.vhd(68[19:45])
    defparam i2425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2424_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_223_0), .O(n2672));   // src/ram.vhd(68[19:45])
    defparam i2424_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1863_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_152_7), .O(n2111));   // src/ram.vhd(68[19:45])
    defparam i1863_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1862_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_152_6), .O(n2110));   // src/ram.vhd(68[19:45])
    defparam i1862_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1861_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_152_5), .O(n2109));   // src/ram.vhd(68[19:45])
    defparam i1861_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1860_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_152_4), .O(n2108));   // src/ram.vhd(68[19:45])
    defparam i1860_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1463_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_102_7), .O(n1711));   // src/ram.vhd(68[19:45])
    defparam i1463_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1462_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_102_6), .O(n1710));   // src/ram.vhd(68[19:45])
    defparam i1462_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1300_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_82_4), .O(n1548));   // src/ram.vhd(68[19:45])
    defparam i1300_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1859_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_152_3), .O(n2107));   // src/ram.vhd(68[19:45])
    defparam i1859_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1461_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_102_5), .O(n1709));   // src/ram.vhd(68[19:45])
    defparam i1461_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1460_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_102_4), .O(n1708));   // src/ram.vhd(68[19:45])
    defparam i1460_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1858_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_152_2), .O(n2106));   // src/ram.vhd(68[19:45])
    defparam i1858_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1459_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_102_3), .O(n1707));   // src/ram.vhd(68[19:45])
    defparam i1459_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1857_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_152_1), .O(n2105));   // src/ram.vhd(68[19:45])
    defparam i1857_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1856_3_lut_4_lut (.I0(n184_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_152_0), .O(n2104));   // src/ram.vhd(68[19:45])
    defparam i1856_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1458_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_102_2), .O(n1706));   // src/ram.vhd(68[19:45])
    defparam i1458_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i35_2_lut (.I0(n19), .I1(port_id[3]), .I2(wea[0]), 
            .I3(wea[0]), .O(n35));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i35_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1457_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_102_1), .O(n1705));   // src/ram.vhd(68[19:45])
    defparam i1457_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1456_3_lut_4_lut (.I0(n211), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_102_0), .O(n1704));   // src/ram.vhd(68[19:45])
    defparam i1456_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2423_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_222_7), .O(n2671));   // src/ram.vhd(68[19:45])
    defparam i2423_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2422_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_222_6), .O(n2670));   // src/ram.vhd(68[19:45])
    defparam i2422_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2421_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_222_5), .O(n2669));   // src/ram.vhd(68[19:45])
    defparam i2421_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1299_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_82_3), .O(n1547));   // src/ram.vhd(68[19:45])
    defparam i1299_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8931_3_lut (.I0(ram_s_208_4), .I1(ram_s_209_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9990));
    defparam i8931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8932_3_lut (.I0(ram_s_210_4), .I1(ram_s_211_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9991));
    defparam i8932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1855_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_151_7), .O(n2103));   // src/ram.vhd(68[19:45])
    defparam i1855_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8941_3_lut (.I0(ram_s_214_4), .I1(ram_s_215_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10000));
    defparam i8941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8940_3_lut (.I0(ram_s_212_4), .I1(ram_s_213_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9999));
    defparam i8940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2420_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_222_4), .O(n2668));   // src/ram.vhd(68[19:45])
    defparam i2420_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1854_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_151_6), .O(n2102));   // src/ram.vhd(68[19:45])
    defparam i1854_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2419_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_222_3), .O(n2667));   // src/ram.vhd(68[19:45])
    defparam i2419_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i25_2_lut (.I0(n18), .I1(port_id[3]), .I2(wea[0]), 
            .I3(wea[0]), .O(n25));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i25_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1853_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_151_5), .O(n2101));   // src/ram.vhd(68[19:45])
    defparam i1853_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1852_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_151_4), .O(n2100));   // src/ram.vhd(68[19:45])
    defparam i1852_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2418_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_222_2), .O(n2666));   // src/ram.vhd(68[19:45])
    defparam i2418_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2417_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_222_1), .O(n2665));   // src/ram.vhd(68[19:45])
    defparam i2417_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2416_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_222_0), .O(n2664));   // src/ram.vhd(68[19:45])
    defparam i2416_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i154_2_lut (.I0(n90_c), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n154));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i154_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2415_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_221_7), .O(n2663));   // src/ram.vhd(68[19:45])
    defparam i2415_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1851_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_151_3), .O(n2099));   // src/ram.vhd(68[19:45])
    defparam i1851_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8001_3_lut (.I0(ram_s_152_5), .I1(ram_s_153_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9060));
    defparam i8001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8002_3_lut (.I0(ram_s_154_5), .I1(ram_s_155_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9061));
    defparam i8002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1850_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_151_2), .O(n2098));   // src/ram.vhd(68[19:45])
    defparam i1850_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2414_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_221_6), .O(n2662));   // src/ram.vhd(68[19:45])
    defparam i2414_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1849_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_151_1), .O(n2097));   // src/ram.vhd(68[19:45])
    defparam i1849_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1848_3_lut_4_lut (.I0(n182_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_151_0), .O(n2096));   // src/ram.vhd(68[19:45])
    defparam i1848_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8077_3_lut (.I0(ram_s_158_5), .I1(ram_s_159_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9136));
    defparam i8077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8076_3_lut (.I0(ram_s_156_5), .I1(ram_s_157_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9135));
    defparam i8076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2413_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_221_5), .O(n2661));   // src/ram.vhd(68[19:45])
    defparam i2413_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2412_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_221_4), .O(n2660));   // src/ram.vhd(68[19:45])
    defparam i2412_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2411_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_221_3), .O(n2659));   // src/ram.vhd(68[19:45])
    defparam i2411_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2410_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_221_2), .O(n2658));   // src/ram.vhd(68[19:45])
    defparam i2410_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2409_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_221_1), .O(n2657));   // src/ram.vhd(68[19:45])
    defparam i2409_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1847_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_150_7), .O(n2095));   // src/ram.vhd(68[19:45])
    defparam i1847_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8067_3_lut (.I0(ram_s_160_0), .I1(ram_s_161_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9126));
    defparam i8067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8068_3_lut (.I0(ram_s_162_0), .I1(ram_s_163_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9127));
    defparam i8068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1846_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_150_6), .O(n2094));   // src/ram.vhd(68[19:45])
    defparam i1846_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1845_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_150_5), .O(n2093));   // src/ram.vhd(68[19:45])
    defparam i1845_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8083_3_lut (.I0(ram_s_166_0), .I1(ram_s_167_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9142));
    defparam i8083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8082_3_lut (.I0(ram_s_164_0), .I1(ram_s_165_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9141));
    defparam i8082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2408_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_221_0), .O(n2656));   // src/ram.vhd(68[19:45])
    defparam i2408_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1844_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_150_4), .O(n2092));   // src/ram.vhd(68[19:45])
    defparam i1844_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8754_3_lut (.I0(ram_s_88_7), .I1(ram_s_89_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9813));
    defparam i8754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8755_3_lut (.I0(ram_s_90_7), .I1(ram_s_91_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9814));
    defparam i8755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1843_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_150_3), .O(n2091));   // src/ram.vhd(68[19:45])
    defparam i1843_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8797_3_lut (.I0(ram_s_94_7), .I1(ram_s_95_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9856));
    defparam i8797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8796_3_lut (.I0(ram_s_92_7), .I1(ram_s_93_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9855));
    defparam i8796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1842_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_150_2), .O(n2090));   // src/ram.vhd(68[19:45])
    defparam i1842_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1841_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_150_1), .O(n2089));   // src/ram.vhd(68[19:45])
    defparam i1841_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i194_2_lut_3_lut (.I0(n65_adj_860), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n194_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i194_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1840_3_lut_4_lut (.I0(n180), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_150_0), .O(n2088));   // src/ram.vhd(68[19:45])
    defparam i1840_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i193_2_lut_3_lut (.I0(n65_adj_860), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n193_adj_859));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i193_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1455_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_101_7), .O(n1703));   // src/ram.vhd(68[19:45])
    defparam i1455_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1454_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_101_6), .O(n1702));   // src/ram.vhd(68[19:45])
    defparam i1454_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1298_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_82_2), .O(n1546));   // src/ram.vhd(68[19:45])
    defparam i1298_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1297_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_82_1), .O(n1545));   // src/ram.vhd(68[19:45])
    defparam i1297_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1296_3_lut_4_lut (.I0(n171), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_82_0), .O(n1544));   // src/ram.vhd(68[19:45])
    defparam i1296_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1453_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_101_5), .O(n1701));   // src/ram.vhd(68[19:45])
    defparam i1453_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1287_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_80_7), .O(n1535));   // src/ram.vhd(68[19:45])
    defparam i1287_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1452_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_101_4), .O(n1700));   // src/ram.vhd(68[19:45])
    defparam i1452_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1451_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_101_3), .O(n1699));   // src/ram.vhd(68[19:45])
    defparam i1451_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1450_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_101_2), .O(n1698));   // src/ram.vhd(68[19:45])
    defparam i1450_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1449_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_101_1), .O(n1697));   // src/ram.vhd(68[19:45])
    defparam i1449_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1448_3_lut_4_lut (.I0(n209), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_101_0), .O(n1696));   // src/ram.vhd(68[19:45])
    defparam i1448_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1839_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_149_7), .O(n2087));   // src/ram.vhd(68[19:45])
    defparam i1839_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2407_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_220_7), .O(n2655));   // src/ram.vhd(68[19:45])
    defparam i2407_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1838_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_149_6), .O(n2086));   // src/ram.vhd(68[19:45])
    defparam i1838_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1837_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_149_5), .O(n2085));   // src/ram.vhd(68[19:45])
    defparam i1837_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2406_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_220_6), .O(n2654));   // src/ram.vhd(68[19:45])
    defparam i2406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2405_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_220_5), .O(n2653));   // src/ram.vhd(68[19:45])
    defparam i2405_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1836_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_149_4), .O(n2084));   // src/ram.vhd(68[19:45])
    defparam i1836_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1835_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_149_3), .O(n2083));   // src/ram.vhd(68[19:45])
    defparam i1835_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1834_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_149_2), .O(n2082));   // src/ram.vhd(68[19:45])
    defparam i1834_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2404_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_220_4), .O(n2652));   // src/ram.vhd(68[19:45])
    defparam i2404_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2403_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_220_3), .O(n2651));   // src/ram.vhd(68[19:45])
    defparam i2403_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1833_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_149_1), .O(n2081));   // src/ram.vhd(68[19:45])
    defparam i1833_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1832_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_149_0), .O(n2080));   // src/ram.vhd(68[19:45])
    defparam i1832_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1286_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_80_6), .O(n1534));   // src/ram.vhd(68[19:45])
    defparam i1286_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1285_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_80_5), .O(n1533));   // src/ram.vhd(68[19:45])
    defparam i1285_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2402_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_220_2), .O(n2650));   // src/ram.vhd(68[19:45])
    defparam i2402_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2401_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_220_1), .O(n2649));   // src/ram.vhd(68[19:45])
    defparam i2401_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8103_3_lut (.I0(ram_s_176_0), .I1(ram_s_177_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9162));
    defparam i8103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8104_3_lut (.I0(ram_s_178_0), .I1(ram_s_179_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9163));
    defparam i8104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8113_3_lut (.I0(ram_s_182_0), .I1(ram_s_183_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9172));
    defparam i8113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8112_3_lut (.I0(ram_s_180_0), .I1(ram_s_181_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9171));
    defparam i8112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1831_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_148_7), .O(n2079));   // src/ram.vhd(68[19:45])
    defparam i1831_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2400_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_220_0), .O(n2648));   // src/ram.vhd(68[19:45])
    defparam i2400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1830_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_148_6), .O(n2078));   // src/ram.vhd(68[19:45])
    defparam i1830_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1829_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_148_5), .O(n2077));   // src/ram.vhd(68[19:45])
    defparam i1829_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8193_3_lut (.I0(ram_s_56_6), .I1(ram_s_57_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9252));
    defparam i8193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8194_3_lut (.I0(ram_s_58_6), .I1(ram_s_59_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9253));
    defparam i8194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i192_2_lut_3_lut (.I0(n63_adj_862), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n192_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i192_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i191_2_lut_3_lut (.I0(n63_adj_862), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n191_adj_861));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i191_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1828_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_148_4), .O(n2076));   // src/ram.vhd(68[19:45])
    defparam i1828_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1827_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_148_3), .O(n2075));   // src/ram.vhd(68[19:45])
    defparam i1827_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1826_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_148_2), .O(n2074));   // src/ram.vhd(68[19:45])
    defparam i1826_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8206_3_lut (.I0(ram_s_62_6), .I1(ram_s_63_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9265));
    defparam i8206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1447_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_100_7), .O(n1695));   // src/ram.vhd(68[19:45])
    defparam i1447_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8205_3_lut (.I0(ram_s_60_6), .I1(ram_s_61_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9264));
    defparam i8205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1825_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_148_1), .O(n2073));   // src/ram.vhd(68[19:45])
    defparam i1825_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8136_3_lut (.I0(ram_s_192_0), .I1(ram_s_193_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9195));
    defparam i8136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1824_3_lut_4_lut (.I0(n176_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_148_0), .O(n2072));   // src/ram.vhd(68[19:45])
    defparam i1824_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1823_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_147_7), .O(n2071));   // src/ram.vhd(68[19:45])
    defparam i1823_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1822_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_147_6), .O(n2070));   // src/ram.vhd(68[19:45])
    defparam i1822_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8137_3_lut (.I0(ram_s_194_0), .I1(ram_s_195_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9196));
    defparam i8137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8149_3_lut (.I0(ram_s_198_0), .I1(ram_s_199_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9208));
    defparam i8149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1821_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_147_5), .O(n2069));   // src/ram.vhd(68[19:45])
    defparam i1821_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8148_3_lut (.I0(ram_s_196_0), .I1(ram_s_197_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9207));
    defparam i8148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1820_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_147_4), .O(n2068));   // src/ram.vhd(68[19:45])
    defparam i1820_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1819_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_147_3), .O(n2067));   // src/ram.vhd(68[19:45])
    defparam i1819_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1818_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_147_2), .O(n2066));   // src/ram.vhd(68[19:45])
    defparam i1818_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1817_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_147_1), .O(n2065));   // src/ram.vhd(68[19:45])
    defparam i1817_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1446_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_100_6), .O(n1694));   // src/ram.vhd(68[19:45])
    defparam i1446_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1816_3_lut_4_lut (.I0(n174), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_147_0), .O(n2064));   // src/ram.vhd(68[19:45])
    defparam i1816_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1445_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_100_5), .O(n1693));   // src/ram.vhd(68[19:45])
    defparam i1445_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1444_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_100_4), .O(n1692));   // src/ram.vhd(68[19:45])
    defparam i1444_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1815_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_146_7), .O(n2063));   // src/ram.vhd(68[19:45])
    defparam i1815_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1284_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_80_4), .O(n1532));   // src/ram.vhd(68[19:45])
    defparam i1284_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1814_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_146_6), .O(n2062));   // src/ram.vhd(68[19:45])
    defparam i1814_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8172_3_lut (.I0(ram_s_208_0), .I1(ram_s_209_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9231));
    defparam i8172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8173_3_lut (.I0(ram_s_210_0), .I1(ram_s_211_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9232));
    defparam i8173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1813_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_146_5), .O(n2061));   // src/ram.vhd(68[19:45])
    defparam i1813_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1812_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_146_4), .O(n2060));   // src/ram.vhd(68[19:45])
    defparam i1812_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1811_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_146_3), .O(n2059));   // src/ram.vhd(68[19:45])
    defparam i1811_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1810_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_146_2), .O(n2058));   // src/ram.vhd(68[19:45])
    defparam i1810_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1443_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_100_3), .O(n1691));   // src/ram.vhd(68[19:45])
    defparam i1443_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i473_474 (.Q(ram_s_19_1), .C(CLK_3P3_MHZ_c), .D(n914));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1442_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_100_2), .O(n1690));   // src/ram.vhd(68[19:45])
    defparam i1442_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1809_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_146_1), .O(n2057));   // src/ram.vhd(68[19:45])
    defparam i1809_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1441_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_100_1), .O(n1689));   // src/ram.vhd(68[19:45])
    defparam i1441_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1808_3_lut_4_lut (.I0(n172), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_146_0), .O(n2056));   // src/ram.vhd(68[19:45])
    defparam i1808_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1440_3_lut_4_lut (.I0(n207), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_100_0), .O(n1688));   // src/ram.vhd(68[19:45])
    defparam i1440_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11483 (.I0(port_id[0]), .I1(ram_s_122_7), 
            .I2(ram_s_123_7), .I3(port_id[1]), .O(n12821));
    defparam port_id_0__bdd_4_lut_11483.LUT_INIT = 16'he4aa;
    SB_LUT4 n12821_bdd_4_lut (.I0(n12821), .I1(ram_s_121_7), .I2(ram_s_120_7), 
            .I3(port_id[1]), .O(n10088));
    defparam n12821_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1807_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_145_7), .O(n2055));   // src/ram.vhd(68[19:45])
    defparam i1807_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1806_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_145_6), .O(n2054));   // src/ram.vhd(68[19:45])
    defparam i1806_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1805_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_145_5), .O(n2053));   // src/ram.vhd(68[19:45])
    defparam i1805_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1804_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_145_4), .O(n2052));   // src/ram.vhd(68[19:45])
    defparam i1804_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1803_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_145_3), .O(n2051));   // src/ram.vhd(68[19:45])
    defparam i1803_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1802_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_145_2), .O(n2050));   // src/ram.vhd(68[19:45])
    defparam i1802_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1801_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_145_1), .O(n2049));   // src/ram.vhd(68[19:45])
    defparam i1801_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1800_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_145_0), .O(n2048));   // src/ram.vhd(68[19:45])
    defparam i1800_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1799_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_144_7), .O(n2047));   // src/ram.vhd(68[19:45])
    defparam i1799_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1798_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_144_6), .O(n2046));   // src/ram.vhd(68[19:45])
    defparam i1798_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1797_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_144_5), .O(n2045));   // src/ram.vhd(68[19:45])
    defparam i1797_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1796_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_144_4), .O(n2044));   // src/ram.vhd(68[19:45])
    defparam i1796_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1795_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_144_3), .O(n2043));   // src/ram.vhd(68[19:45])
    defparam i1795_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1794_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_144_2), .O(n2042));   // src/ram.vhd(68[19:45])
    defparam i1794_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1793_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_144_1), .O(n2041));   // src/ram.vhd(68[19:45])
    defparam i1793_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1792_3_lut_4_lut (.I0(n168), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_144_0), .O(n2040));   // src/ram.vhd(68[19:45])
    defparam i1792_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1791_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_143_7), .O(n2039));   // src/ram.vhd(68[19:45])
    defparam i1791_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1790_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_143_6), .O(n2038));   // src/ram.vhd(68[19:45])
    defparam i1790_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1789_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_143_5), .O(n2037));   // src/ram.vhd(68[19:45])
    defparam i1789_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1788_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_143_4), .O(n2036));   // src/ram.vhd(68[19:45])
    defparam i1788_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1787_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_143_3), .O(n2035));   // src/ram.vhd(68[19:45])
    defparam i1787_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1786_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_143_2), .O(n2034));   // src/ram.vhd(68[19:45])
    defparam i1786_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1785_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_143_1), .O(n2033));   // src/ram.vhd(68[19:45])
    defparam i1785_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1784_3_lut_4_lut (.I0(n166), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_143_0), .O(n2032));   // src/ram.vhd(68[19:45])
    defparam i1784_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i649_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_9_6), .O(n897));   // src/ram.vhd(68[19:45])
    defparam i649_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i734_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_9_5), .O(n982));   // src/ram.vhd(68[19:45])
    defparam i734_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i751_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_9_0), .O(n999));   // src/ram.vhd(68[19:45])
    defparam i751_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i733_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_9_2), .O(n981));   // src/ram.vhd(68[19:45])
    defparam i733_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i743_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_9_4), .O(n991));   // src/ram.vhd(68[19:45])
    defparam i743_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i752_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_9_3), .O(n1000));   // src/ram.vhd(68[19:45])
    defparam i752_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i680_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_9_7), .O(n928));   // src/ram.vhd(68[19:45])
    defparam i680_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i742_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_9_1), .O(n990));   // src/ram.vhd(68[19:45])
    defparam i742_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i217_2_lut_3_lut_4_lut (.I0(n25), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n217_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i217_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i218_2_lut_3_lut_4_lut (.I0(n25), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n218_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i218_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 EnabledDecoder_2_i290_2_lut_3_lut (.I0(n98), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n244));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i290_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i289_2_lut_3_lut (.I0(n98), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n116));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i289_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i21_2_lut_3_lut_4_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[2]), .I3(port_id[1]), .O(n21));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i21_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i22_2_lut_3_lut_4_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[2]), .I3(port_id[1]), .O(n22));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i22_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 EnabledDecoder_2_i291_2_lut_3_lut (.I0(n100), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n115));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i291_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i292_2_lut_3_lut (.I0(n100), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n243));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i292_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i288_2_lut_3_lut (.I0(n96_adj_864), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n245));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i288_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i287_2_lut_3_lut (.I0(n96_adj_864), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n117));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i287_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i227_2_lut_3_lut_4_lut (.I0(n35), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n227));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i227_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i228_2_lut_3_lut_4_lut (.I0(n35), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n228));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i228_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i644_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_21_3), .O(n892));   // src/ram.vhd(68[19:45])
    defparam i644_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i815_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_21_7), .O(n1063));   // src/ram.vhd(68[19:45])
    defparam i815_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i657_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_21_2), .O(n905));   // src/ram.vhd(68[19:45])
    defparam i657_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i664_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_21_1), .O(n912));   // src/ram.vhd(68[19:45])
    defparam i664_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i667_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_21_0), .O(n915));   // src/ram.vhd(68[19:45])
    defparam i667_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i808_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_21_4), .O(n1056));   // src/ram.vhd(68[19:45])
    defparam i808_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i813_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_21_5), .O(n1061));   // src/ram.vhd(68[19:45])
    defparam i813_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i814_3_lut_4_lut (.I0(n178), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_21_6), .O(n1062));   // src/ram.vhd(68[19:45])
    defparam i814_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i177_2_lut_3_lut (.I0(n49), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n177));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i177_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i178_2_lut_3_lut (.I0(n49), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n178));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i178_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i49_2_lut_3_lut (.I0(n17), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n49));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i49_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i81_2_lut_3_lut_4_lut (.I0(n17), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n81));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i81_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i82_2_lut_3_lut_4_lut (.I0(n17), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n82_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i82_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i286_2_lut_3_lut (.I0(n94_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n246));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i286_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i285_2_lut_3_lut (.I0(n94_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n118));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i285_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i643_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_17_0), .O(n891));   // src/ram.vhd(68[19:45])
    defparam i643_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i672_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_17_7), .O(n920));   // src/ram.vhd(68[19:45])
    defparam i672_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i791_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_17_6), .O(n1039));   // src/ram.vhd(68[19:45])
    defparam i791_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i637_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_17_5), .O(n885));   // src/ram.vhd(68[19:45])
    defparam i637_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i639_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_17_4), .O(n887));   // src/ram.vhd(68[19:45])
    defparam i639_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i640_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_17_3), .O(n888));   // src/ram.vhd(68[19:45])
    defparam i640_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i641_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_17_2), .O(n889));   // src/ram.vhd(68[19:45])
    defparam i641_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i642_3_lut_4_lut (.I0(n170), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_17_1), .O(n890));   // src/ram.vhd(68[19:45])
    defparam i642_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i170_2_lut_3_lut (.I0(n41), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n170));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i170_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i425_2_lut_3_lut_4_lut (.I0(n41), .I1(port_id[5]), 
            .I2(port_id[7]), .I3(port_id[6]), .O(n48));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i425_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i426_2_lut_3_lut_4_lut (.I0(n41), .I1(port_id[5]), 
            .I2(port_id[7]), .I3(port_id[6]), .O(n176));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i426_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1751_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_138_7), .O(n1999));   // src/ram.vhd(68[19:45])
    defparam i1751_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1750_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_138_6), .O(n1998));   // src/ram.vhd(68[19:45])
    defparam i1750_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1749_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_138_5), .O(n1997));   // src/ram.vhd(68[19:45])
    defparam i1749_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1748_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_138_4), .O(n1996));   // src/ram.vhd(68[19:45])
    defparam i1748_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1747_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_138_3), .O(n1995));   // src/ram.vhd(68[19:45])
    defparam i1747_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1746_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_138_2), .O(n1994));   // src/ram.vhd(68[19:45])
    defparam i1746_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1745_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_138_1), .O(n1993));   // src/ram.vhd(68[19:45])
    defparam i1745_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1744_3_lut_4_lut (.I0(n156), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_138_0), .O(n1992));   // src/ram.vhd(68[19:45])
    defparam i1744_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i41_2_lut_3_lut (.I0(n18), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n41));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i41_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i73_2_lut_3_lut_4_lut (.I0(n18), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n73));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i73_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i74_2_lut_3_lut_4_lut (.I0(n18), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n74));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i74_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1743_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_137_7), .O(n1991));   // src/ram.vhd(68[19:45])
    defparam i1743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1742_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_137_6), .O(n1990));   // src/ram.vhd(68[19:45])
    defparam i1742_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1741_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_137_5), .O(n1989));   // src/ram.vhd(68[19:45])
    defparam i1741_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1740_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_137_4), .O(n1988));   // src/ram.vhd(68[19:45])
    defparam i1740_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1739_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_137_3), .O(n1987));   // src/ram.vhd(68[19:45])
    defparam i1739_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1738_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_137_2), .O(n1986));   // src/ram.vhd(68[19:45])
    defparam i1738_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1737_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_137_1), .O(n1985));   // src/ram.vhd(68[19:45])
    defparam i1737_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1736_3_lut_4_lut (.I0(n154), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_137_0), .O(n1984));   // src/ram.vhd(68[19:45])
    defparam i1736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i280_2_lut_3_lut (.I0(n88), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n249));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i280_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i279_2_lut_3_lut (.I0(n88), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n121));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i279_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i278_2_lut_3_lut (.I0(n86_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n250));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i278_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i277_2_lut_3_lut (.I0(n86_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n122));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i277_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i276_2_lut_3_lut (.I0(n84_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n251));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i276_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i275_2_lut_3_lut (.I0(n84_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n123));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i275_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i274_2_lut_3_lut (.I0(n82_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n252));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i274_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i273_2_lut_3_lut (.I0(n82_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n124));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i273_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i272_2_lut_3_lut (.I0(n80), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n253));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i272_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i271_2_lut_3_lut (.I0(n80), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n125));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i271_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i270_2_lut_3_lut (.I0(n78), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n254));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i270_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i269_2_lut_3_lut (.I0(n78), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n126));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i269_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i268_2_lut_3_lut (.I0(n76), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n255));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i268_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i267_2_lut_3_lut (.I0(n76), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n127));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i267_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i266_2_lut_3_lut (.I0(n74), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n256));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i266_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i265_2_lut_3_lut (.I0(n74), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n128));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i265_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2687_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_255_7), .O(n2935));   // src/ram.vhd(68[19:45])
    defparam i2687_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2686_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_255_6), .O(n2934));   // src/ram.vhd(68[19:45])
    defparam i2686_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2685_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_255_5), .O(n2933));   // src/ram.vhd(68[19:45])
    defparam i2685_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2684_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_255_4), .O(n2932));   // src/ram.vhd(68[19:45])
    defparam i2684_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2683_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_255_3), .O(n2931));   // src/ram.vhd(68[19:45])
    defparam i2683_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2682_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_255_2), .O(n2930));   // src/ram.vhd(68[19:45])
    defparam i2682_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2681_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_255_1), .O(n2929));   // src/ram.vhd(68[19:45])
    defparam i2681_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2680_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_255_0), .O(n2928));   // src/ram.vhd(68[19:45])
    defparam i2680_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i197_2_lut_3_lut_4_lut (.I0(n37), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n197));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i197_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i198_2_lut_3_lut_4_lut (.I0(n37), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n198));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i198_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i264_2_lut_3_lut (.I0(n72_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n257));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i264_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i263_2_lut_3_lut (.I0(n72_c), .I1(port_id[6]), 
            .I2(port_id[7]), .I3(wea[0]), .O(n129));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i263_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2679_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_254_7), .O(n2927));   // src/ram.vhd(68[19:45])
    defparam i2679_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2678_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_254_6), .O(n2926));   // src/ram.vhd(68[19:45])
    defparam i2678_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2677_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_254_5), .O(n2925));   // src/ram.vhd(68[19:45])
    defparam i2677_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2676_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_254_4), .O(n2924));   // src/ram.vhd(68[19:45])
    defparam i2676_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2675_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_254_3), .O(n2923));   // src/ram.vhd(68[19:45])
    defparam i2675_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2674_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_254_2), .O(n2922));   // src/ram.vhd(68[19:45])
    defparam i2674_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2673_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_254_1), .O(n2921));   // src/ram.vhd(68[19:45])
    defparam i2673_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2672_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_254_0), .O(n2920));   // src/ram.vhd(68[19:45])
    defparam i2672_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i195_2_lut_3_lut_4_lut (.I0(n35), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n195_adj_858));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i195_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i196_2_lut_3_lut_4_lut (.I0(n35), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n196));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i196_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i2671_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_253_7), .O(n2919));   // src/ram.vhd(68[19:45])
    defparam i2671_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2670_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_253_6), .O(n2918));   // src/ram.vhd(68[19:45])
    defparam i2670_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2669_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_253_5), .O(n2917));   // src/ram.vhd(68[19:45])
    defparam i2669_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2668_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_253_4), .O(n2916));   // src/ram.vhd(68[19:45])
    defparam i2668_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2667_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_253_3), .O(n2915));   // src/ram.vhd(68[19:45])
    defparam i2667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2666_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_253_2), .O(n2914));   // src/ram.vhd(68[19:45])
    defparam i2666_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2665_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_253_1), .O(n2913));   // src/ram.vhd(68[19:45])
    defparam i2665_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2664_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_253_0), .O(n2912));   // src/ram.vhd(68[19:45])
    defparam i2664_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i258_2_lut_3_lut (.I0(n65_adj_860), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n258));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i258_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i257_2_lut_3_lut (.I0(n65_adj_860), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n257_adj_873));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i257_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1663_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_127_7), .O(n1911));   // src/ram.vhd(68[19:45])
    defparam i1663_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1662_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_127_6), .O(n1910));   // src/ram.vhd(68[19:45])
    defparam i1662_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1661_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_127_5), .O(n1909));   // src/ram.vhd(68[19:45])
    defparam i1661_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1660_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_127_4), .O(n1908));   // src/ram.vhd(68[19:45])
    defparam i1660_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1659_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_127_3), .O(n1907));   // src/ram.vhd(68[19:45])
    defparam i1659_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1658_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_127_2), .O(n1906));   // src/ram.vhd(68[19:45])
    defparam i1658_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1657_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_127_1), .O(n1905));   // src/ram.vhd(68[19:45])
    defparam i1657_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1656_3_lut_4_lut (.I0(n261), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_127_0), .O(n1904));   // src/ram.vhd(68[19:45])
    defparam i1656_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i65_2_lut_3_lut (.I0(n17), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n65_adj_860));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i65_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i97_2_lut_3_lut_4_lut (.I0(n17), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n97_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i97_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i98_2_lut_3_lut_4_lut (.I0(n17), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n98));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i98_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i2663_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_252_7), .O(n2911));   // src/ram.vhd(68[19:45])
    defparam i2663_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2662_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_252_6), .O(n2910));   // src/ram.vhd(68[19:45])
    defparam i2662_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2661_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_252_5), .O(n2909));   // src/ram.vhd(68[19:45])
    defparam i2661_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2660_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_252_4), .O(n2908));   // src/ram.vhd(68[19:45])
    defparam i2660_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2659_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_252_3), .O(n2907));   // src/ram.vhd(68[19:45])
    defparam i2659_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2658_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_252_2), .O(n2906));   // src/ram.vhd(68[19:45])
    defparam i2658_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2657_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_252_1), .O(n2905));   // src/ram.vhd(68[19:45])
    defparam i2657_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2656_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_252_0), .O(n2904));   // src/ram.vhd(68[19:45])
    defparam i2656_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i256_2_lut_3_lut (.I0(n63_adj_862), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n256_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i256_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i255_2_lut_3_lut (.I0(n63_adj_862), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n255_adj_874));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i255_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i63_2_lut_3_lut (.I0(n15), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n63_adj_862));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i63_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i95_2_lut_3_lut_4_lut (.I0(n15), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n95_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i95_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i96_2_lut_3_lut_4_lut (.I0(n15), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n96_adj_864));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i96_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1655_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_126_7), .O(n1903));   // src/ram.vhd(68[19:45])
    defparam i1655_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1654_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_126_6), .O(n1902));   // src/ram.vhd(68[19:45])
    defparam i1654_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1653_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_126_5), .O(n1901));   // src/ram.vhd(68[19:45])
    defparam i1653_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1652_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_126_4), .O(n1900));   // src/ram.vhd(68[19:45])
    defparam i1652_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1651_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_126_3), .O(n1899));   // src/ram.vhd(68[19:45])
    defparam i1651_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1650_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_126_2), .O(n1898));   // src/ram.vhd(68[19:45])
    defparam i1650_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1649_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_126_1), .O(n1897));   // src/ram.vhd(68[19:45])
    defparam i1649_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1648_3_lut_4_lut (.I0(n259), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_126_0), .O(n1896));   // src/ram.vhd(68[19:45])
    defparam i1648_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2655_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_251_7), .O(n2903));   // src/ram.vhd(68[19:45])
    defparam i2655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2654_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_251_6), .O(n2902));   // src/ram.vhd(68[19:45])
    defparam i2654_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2653_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_251_5), .O(n2901));   // src/ram.vhd(68[19:45])
    defparam i2653_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2652_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_251_4), .O(n2900));   // src/ram.vhd(68[19:45])
    defparam i2652_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2651_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_251_3), .O(n2899));   // src/ram.vhd(68[19:45])
    defparam i2651_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2650_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_251_2), .O(n2898));   // src/ram.vhd(68[19:45])
    defparam i2650_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2649_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_251_1), .O(n2897));   // src/ram.vhd(68[19:45])
    defparam i2649_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2648_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_251_0), .O(n2896));   // src/ram.vhd(68[19:45])
    defparam i2648_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i254_2_lut_3_lut (.I0(n61_adj_876), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n254_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i254_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i253_2_lut_3_lut (.I0(n61_adj_876), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n253_adj_875));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i253_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i61_2_lut_3_lut (.I0(n22), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n61_adj_876));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i61_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i93_2_lut_3_lut_4_lut (.I0(n22), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n93_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i93_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i94_2_lut_3_lut_4_lut (.I0(n22), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n94_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i94_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1647_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_125_7), .O(n1895));   // src/ram.vhd(68[19:45])
    defparam i1647_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1646_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_125_6), .O(n1894));   // src/ram.vhd(68[19:45])
    defparam i1646_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1645_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_125_5), .O(n1893));   // src/ram.vhd(68[19:45])
    defparam i1645_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1644_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_125_4), .O(n1892));   // src/ram.vhd(68[19:45])
    defparam i1644_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1643_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_125_3), .O(n1891));   // src/ram.vhd(68[19:45])
    defparam i1643_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1642_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_125_2), .O(n1890));   // src/ram.vhd(68[19:45])
    defparam i1642_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1641_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_125_1), .O(n1889));   // src/ram.vhd(68[19:45])
    defparam i1641_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1640_3_lut_4_lut (.I0(n257_adj_873), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_125_0), .O(n1888));   // src/ram.vhd(68[19:45])
    defparam i1640_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2647_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_250_7), .O(n2895));   // src/ram.vhd(68[19:45])
    defparam i2647_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2646_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_250_6), .O(n2894));   // src/ram.vhd(68[19:45])
    defparam i2646_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2645_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_250_5), .O(n2893));   // src/ram.vhd(68[19:45])
    defparam i2645_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2644_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_250_4), .O(n2892));   // src/ram.vhd(68[19:45])
    defparam i2644_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2643_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_250_3), .O(n2891));   // src/ram.vhd(68[19:45])
    defparam i2643_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2642_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_250_2), .O(n2890));   // src/ram.vhd(68[19:45])
    defparam i2642_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2641_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_250_1), .O(n2889));   // src/ram.vhd(68[19:45])
    defparam i2641_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2640_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_250_0), .O(n2888));   // src/ram.vhd(68[19:45])
    defparam i2640_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i187_2_lut_3_lut_4_lut (.I0(n27), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n187_adj_877));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i187_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i188_2_lut_3_lut_4_lut (.I0(n27), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n188_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i188_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i2639_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_249_7), .O(n2887));   // src/ram.vhd(68[19:45])
    defparam i2639_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2638_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_249_6), .O(n2886));   // src/ram.vhd(68[19:45])
    defparam i2638_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2637_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_249_5), .O(n2885));   // src/ram.vhd(68[19:45])
    defparam i2637_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2636_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_249_4), .O(n2884));   // src/ram.vhd(68[19:45])
    defparam i2636_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2635_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_249_3), .O(n2883));   // src/ram.vhd(68[19:45])
    defparam i2635_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2634_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_249_2), .O(n2882));   // src/ram.vhd(68[19:45])
    defparam i2634_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2633_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_249_1), .O(n2881));   // src/ram.vhd(68[19:45])
    defparam i2633_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2632_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_249_0), .O(n2880));   // src/ram.vhd(68[19:45])
    defparam i2632_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1639_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_124_7), .O(n1887));   // src/ram.vhd(68[19:45])
    defparam i1639_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1638_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_124_6), .O(n1886));   // src/ram.vhd(68[19:45])
    defparam i1638_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1637_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_124_5), .O(n1885));   // src/ram.vhd(68[19:45])
    defparam i1637_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1636_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_124_4), .O(n1884));   // src/ram.vhd(68[19:45])
    defparam i1636_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1635_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_124_3), .O(n1883));   // src/ram.vhd(68[19:45])
    defparam i1635_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1634_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_124_2), .O(n1882));   // src/ram.vhd(68[19:45])
    defparam i1634_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1633_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_124_1), .O(n1881));   // src/ram.vhd(68[19:45])
    defparam i1633_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1632_3_lut_4_lut (.I0(n255_adj_874), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_124_0), .O(n1880));   // src/ram.vhd(68[19:45])
    defparam i1632_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i185_2_lut_3_lut_4_lut (.I0(n25), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n185_adj_878));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i185_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i186_2_lut_3_lut_4_lut (.I0(n25), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n186_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i186_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i2631_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_248_7), .O(n2879));   // src/ram.vhd(68[19:45])
    defparam i2631_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2630_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_248_6), .O(n2878));   // src/ram.vhd(68[19:45])
    defparam i2630_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2629_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_248_5), .O(n2877));   // src/ram.vhd(68[19:45])
    defparam i2629_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2628_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_248_4), .O(n2876));   // src/ram.vhd(68[19:45])
    defparam i2628_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2627_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_248_3), .O(n2875));   // src/ram.vhd(68[19:45])
    defparam i2627_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2626_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_248_2), .O(n2874));   // src/ram.vhd(68[19:45])
    defparam i2626_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2625_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_248_1), .O(n2873));   // src/ram.vhd(68[19:45])
    defparam i2625_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2624_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_248_0), .O(n2872));   // src/ram.vhd(68[19:45])
    defparam i2624_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i248_2_lut_3_lut (.I0(n55_adj_879), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n248));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i248_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i247_2_lut_3_lut (.I0(n55_adj_879), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n247));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i247_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i55_2_lut_3_lut (.I0(n16), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n55_adj_879));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i55_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i87_2_lut_3_lut_4_lut (.I0(n16), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n87));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i87_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i88_2_lut_3_lut_4_lut (.I0(n16), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n88));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i88_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1631_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_123_7), .O(n1879));   // src/ram.vhd(68[19:45])
    defparam i1631_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1630_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_123_6), .O(n1878));   // src/ram.vhd(68[19:45])
    defparam i1630_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1629_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_123_5), .O(n1877));   // src/ram.vhd(68[19:45])
    defparam i1629_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1628_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_123_4), .O(n1876));   // src/ram.vhd(68[19:45])
    defparam i1628_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1627_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_123_3), .O(n1875));   // src/ram.vhd(68[19:45])
    defparam i1627_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1626_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_123_2), .O(n1874));   // src/ram.vhd(68[19:45])
    defparam i1626_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1625_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_123_1), .O(n1873));   // src/ram.vhd(68[19:45])
    defparam i1625_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1624_3_lut_4_lut (.I0(n253_adj_875), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_123_0), .O(n1872));   // src/ram.vhd(68[19:45])
    defparam i1624_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2623_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_247_7), .O(n2871));   // src/ram.vhd(68[19:45])
    defparam i2623_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2622_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_247_6), .O(n2870));   // src/ram.vhd(68[19:45])
    defparam i2622_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2621_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_247_5), .O(n2869));   // src/ram.vhd(68[19:45])
    defparam i2621_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2620_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_247_4), .O(n2868));   // src/ram.vhd(68[19:45])
    defparam i2620_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2619_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_247_3), .O(n2867));   // src/ram.vhd(68[19:45])
    defparam i2619_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2618_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_247_2), .O(n2866));   // src/ram.vhd(68[19:45])
    defparam i2618_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2617_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_247_1), .O(n2865));   // src/ram.vhd(68[19:45])
    defparam i2617_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2616_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_247_0), .O(n2864));   // src/ram.vhd(68[19:45])
    defparam i2616_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i246_2_lut_3_lut (.I0(n53), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n246_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i246_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i245_2_lut_3_lut (.I0(n53), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n245_adj_880));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i245_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i53_2_lut_3_lut (.I0(n21), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n53));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i53_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i85_2_lut_3_lut_4_lut (.I0(n21), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n85_adj_845));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i85_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i86_2_lut_3_lut_4_lut (.I0(n21), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n86_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i86_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1623_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_122_7), .O(n1871));   // src/ram.vhd(68[19:45])
    defparam i1623_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1622_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_122_6), .O(n1870));   // src/ram.vhd(68[19:45])
    defparam i1622_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1621_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_122_5), .O(n1869));   // src/ram.vhd(68[19:45])
    defparam i1621_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1620_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_122_4), .O(n1868));   // src/ram.vhd(68[19:45])
    defparam i1620_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1619_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_122_3), .O(n1867));   // src/ram.vhd(68[19:45])
    defparam i1619_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1618_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_122_2), .O(n1866));   // src/ram.vhd(68[19:45])
    defparam i1618_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1617_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_122_1), .O(n1865));   // src/ram.vhd(68[19:45])
    defparam i1617_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1616_3_lut_4_lut (.I0(n251_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_122_0), .O(n1864));   // src/ram.vhd(68[19:45])
    defparam i1616_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2615_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_246_7), .O(n2863));   // src/ram.vhd(68[19:45])
    defparam i2615_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2614_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_246_6), .O(n2862));   // src/ram.vhd(68[19:45])
    defparam i2614_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2613_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_246_5), .O(n2861));   // src/ram.vhd(68[19:45])
    defparam i2613_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2612_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_246_4), .O(n2860));   // src/ram.vhd(68[19:45])
    defparam i2612_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2611_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_246_3), .O(n2859));   // src/ram.vhd(68[19:45])
    defparam i2611_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2610_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_246_2), .O(n2858));   // src/ram.vhd(68[19:45])
    defparam i2610_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2609_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_246_1), .O(n2857));   // src/ram.vhd(68[19:45])
    defparam i2609_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2608_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_246_0), .O(n2856));   // src/ram.vhd(68[19:45])
    defparam i2608_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i244_2_lut_3_lut (.I0(n51), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n244_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i244_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i243_2_lut_3_lut (.I0(n51), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n243_adj_881));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i243_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i51_2_lut_3_lut (.I0(n19), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n51));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i51_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i83_2_lut_3_lut_4_lut (.I0(n19), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n83));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i83_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i84_2_lut_3_lut_4_lut (.I0(n19), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n84_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i84_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1615_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_121_7), .O(n1863));   // src/ram.vhd(68[19:45])
    defparam i1615_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1614_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_121_6), .O(n1862));   // src/ram.vhd(68[19:45])
    defparam i1614_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1613_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_121_5), .O(n1861));   // src/ram.vhd(68[19:45])
    defparam i1613_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1612_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_121_4), .O(n1860));   // src/ram.vhd(68[19:45])
    defparam i1612_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1611_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_121_3), .O(n1859));   // src/ram.vhd(68[19:45])
    defparam i1611_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1610_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_121_2), .O(n1858));   // src/ram.vhd(68[19:45])
    defparam i1610_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1609_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_121_1), .O(n1857));   // src/ram.vhd(68[19:45])
    defparam i1609_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1608_3_lut_4_lut (.I0(n249_c), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_121_0), .O(n1856));   // src/ram.vhd(68[19:45])
    defparam i1608_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2607_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_245_7), .O(n2855));   // src/ram.vhd(68[19:45])
    defparam i2607_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2606_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_245_6), .O(n2854));   // src/ram.vhd(68[19:45])
    defparam i2606_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2605_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_245_5), .O(n2853));   // src/ram.vhd(68[19:45])
    defparam i2605_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2604_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_245_4), .O(n2852));   // src/ram.vhd(68[19:45])
    defparam i2604_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2603_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_245_3), .O(n2851));   // src/ram.vhd(68[19:45])
    defparam i2603_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2602_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_245_2), .O(n2850));   // src/ram.vhd(68[19:45])
    defparam i2602_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2601_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_245_1), .O(n2849));   // src/ram.vhd(68[19:45])
    defparam i2601_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2600_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_245_0), .O(n2848));   // src/ram.vhd(68[19:45])
    defparam i2600_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i242_2_lut_3_lut (.I0(n49), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n242));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i242_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i241_2_lut_3_lut (.I0(n49), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n241));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i241_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2599_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_244_7), .O(n2847));   // src/ram.vhd(68[19:45])
    defparam i2599_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2598_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_244_6), .O(n2846));   // src/ram.vhd(68[19:45])
    defparam i2598_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2597_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_244_5), .O(n2845));   // src/ram.vhd(68[19:45])
    defparam i2597_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2596_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_244_4), .O(n2844));   // src/ram.vhd(68[19:45])
    defparam i2596_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2595_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_244_3), .O(n2843));   // src/ram.vhd(68[19:45])
    defparam i2595_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2594_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_244_2), .O(n2842));   // src/ram.vhd(68[19:45])
    defparam i2594_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2593_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_244_1), .O(n2841));   // src/ram.vhd(68[19:45])
    defparam i2593_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2399_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_219_7), .O(n2647));   // src/ram.vhd(68[19:45])
    defparam i2399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2398_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_219_6), .O(n2646));   // src/ram.vhd(68[19:45])
    defparam i2398_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2397_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_219_5), .O(n2645));   // src/ram.vhd(68[19:45])
    defparam i2397_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2396_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_219_4), .O(n2644));   // src/ram.vhd(68[19:45])
    defparam i2396_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2592_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_244_0), .O(n2840));   // src/ram.vhd(68[19:45])
    defparam i2592_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i240_2_lut_3_lut (.I0(n47), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n240));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i240_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i239_2_lut_3_lut (.I0(n47), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n239));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i239_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut (.I0(n15), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n47));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i47_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i79_2_lut_3_lut_4_lut (.I0(n15), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n79));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i79_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i80_2_lut_3_lut_4_lut (.I0(n15), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n80));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i80_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1607_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_120_7), .O(n1855));   // src/ram.vhd(68[19:45])
    defparam i1607_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1606_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_120_6), .O(n1854));   // src/ram.vhd(68[19:45])
    defparam i1606_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1605_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_120_5), .O(n1853));   // src/ram.vhd(68[19:45])
    defparam i1605_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1604_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_120_4), .O(n1852));   // src/ram.vhd(68[19:45])
    defparam i1604_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1603_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_120_3), .O(n1851));   // src/ram.vhd(68[19:45])
    defparam i1603_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1602_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_120_2), .O(n1850));   // src/ram.vhd(68[19:45])
    defparam i1602_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1601_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_120_1), .O(n1849));   // src/ram.vhd(68[19:45])
    defparam i1601_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1600_3_lut_4_lut (.I0(n247), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_120_0), .O(n1848));   // src/ram.vhd(68[19:45])
    defparam i1600_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2591_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_243_7), .O(n2839));   // src/ram.vhd(68[19:45])
    defparam i2591_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2590_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_243_6), .O(n2838));   // src/ram.vhd(68[19:45])
    defparam i2590_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2589_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_243_5), .O(n2837));   // src/ram.vhd(68[19:45])
    defparam i2589_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2588_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_243_4), .O(n2836));   // src/ram.vhd(68[19:45])
    defparam i2588_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2587_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_243_3), .O(n2835));   // src/ram.vhd(68[19:45])
    defparam i2587_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2586_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_243_2), .O(n2834));   // src/ram.vhd(68[19:45])
    defparam i2586_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2585_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_243_1), .O(n2833));   // src/ram.vhd(68[19:45])
    defparam i2585_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2584_3_lut_4_lut (.I0(n237), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_243_0), .O(n2832));   // src/ram.vhd(68[19:45])
    defparam i2584_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i238_2_lut_3_lut (.I0(n45), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n238));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i238_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i237_2_lut_3_lut (.I0(n45), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n237));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i237_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut (.I0(n22), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n45));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i45_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i77_2_lut_3_lut_4_lut (.I0(n22), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n77));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i77_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i78_2_lut_3_lut_4_lut (.I0(n22), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n78));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i78_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1599_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_119_7), .O(n1847));   // src/ram.vhd(68[19:45])
    defparam i1599_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1598_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_119_6), .O(n1846));   // src/ram.vhd(68[19:45])
    defparam i1598_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1597_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_119_5), .O(n1845));   // src/ram.vhd(68[19:45])
    defparam i1597_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1596_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_119_4), .O(n1844));   // src/ram.vhd(68[19:45])
    defparam i1596_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1595_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_119_3), .O(n1843));   // src/ram.vhd(68[19:45])
    defparam i1595_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1594_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_119_2), .O(n1842));   // src/ram.vhd(68[19:45])
    defparam i1594_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1593_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_119_1), .O(n1841));   // src/ram.vhd(68[19:45])
    defparam i1593_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1592_3_lut_4_lut (.I0(n245_adj_880), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_119_0), .O(n1840));   // src/ram.vhd(68[19:45])
    defparam i1592_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2583_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_242_7), .O(n2831));   // src/ram.vhd(68[19:45])
    defparam i2583_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2582_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_242_6), .O(n2830));   // src/ram.vhd(68[19:45])
    defparam i2582_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2581_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_242_5), .O(n2829));   // src/ram.vhd(68[19:45])
    defparam i2581_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2580_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_242_4), .O(n2828));   // src/ram.vhd(68[19:45])
    defparam i2580_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2579_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_242_3), .O(n2827));   // src/ram.vhd(68[19:45])
    defparam i2579_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2578_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_242_2), .O(n2826));   // src/ram.vhd(68[19:45])
    defparam i2578_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2577_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_242_1), .O(n2825));   // src/ram.vhd(68[19:45])
    defparam i2577_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2576_3_lut_4_lut (.I0(n235), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_242_0), .O(n2824));   // src/ram.vhd(68[19:45])
    defparam i2576_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i236_2_lut_3_lut (.I0(n43), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n236));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i236_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i235_2_lut_3_lut (.I0(n43), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n235));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i235_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i75_2_lut_3_lut_4_lut (.I0(n20), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n75));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i75_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i76_2_lut_3_lut_4_lut (.I0(n20), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n76));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i76_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i2575_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_241_7), .O(n2823));   // src/ram.vhd(68[19:45])
    defparam i2575_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2574_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_241_6), .O(n2822));   // src/ram.vhd(68[19:45])
    defparam i2574_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2573_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_241_5), .O(n2821));   // src/ram.vhd(68[19:45])
    defparam i2573_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2572_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_241_4), .O(n2820));   // src/ram.vhd(68[19:45])
    defparam i2572_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2571_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_241_3), .O(n2819));   // src/ram.vhd(68[19:45])
    defparam i2571_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2570_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_241_2), .O(n2818));   // src/ram.vhd(68[19:45])
    defparam i2570_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2569_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_241_1), .O(n2817));   // src/ram.vhd(68[19:45])
    defparam i2569_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2568_3_lut_4_lut (.I0(n233), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_241_0), .O(n2816));   // src/ram.vhd(68[19:45])
    defparam i2568_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1591_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_118_7), .O(n1839));   // src/ram.vhd(68[19:45])
    defparam i1591_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1590_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_118_6), .O(n1838));   // src/ram.vhd(68[19:45])
    defparam i1590_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1589_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_118_5), .O(n1837));   // src/ram.vhd(68[19:45])
    defparam i1589_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2395_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_219_3), .O(n2643));   // src/ram.vhd(68[19:45])
    defparam i2395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2394_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_219_2), .O(n2642));   // src/ram.vhd(68[19:45])
    defparam i2394_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2393_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_219_1), .O(n2641));   // src/ram.vhd(68[19:45])
    defparam i2393_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2392_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_219_0), .O(n2640));   // src/ram.vhd(68[19:45])
    defparam i2392_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i190_2_lut_3_lut (.I0(n61_adj_876), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n190_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i190_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i189_2_lut_3_lut (.I0(n61_adj_876), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n189_adj_882));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i189_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1439_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_99_7), .O(n1687));   // src/ram.vhd(68[19:45])
    defparam i1439_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1438_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_99_6), .O(n1686));   // src/ram.vhd(68[19:45])
    defparam i1438_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1283_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_80_3), .O(n1531));   // src/ram.vhd(68[19:45])
    defparam i1283_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1282_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_80_2), .O(n1530));   // src/ram.vhd(68[19:45])
    defparam i1282_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1437_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_99_5), .O(n1685));   // src/ram.vhd(68[19:45])
    defparam i1437_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1588_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_118_4), .O(n1836));   // src/ram.vhd(68[19:45])
    defparam i1588_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8182_3_lut (.I0(ram_s_214_0), .I1(ram_s_215_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9241));
    defparam i8182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8181_3_lut (.I0(ram_s_212_0), .I1(ram_s_213_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9240));
    defparam i8181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2297_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_207_1), .O(n2545));   // src/ram.vhd(68[19:45])
    defparam i2297_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1281_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_80_1), .O(n1529));   // src/ram.vhd(68[19:45])
    defparam i1281_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2296_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_207_0), .O(n2544));   // src/ram.vhd(68[19:45])
    defparam i2296_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1436_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_99_4), .O(n1684));   // src/ram.vhd(68[19:45])
    defparam i1436_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1280_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_80_0), .O(n1528));   // src/ram.vhd(68[19:45])
    defparam i1280_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1435_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_99_3), .O(n1683));   // src/ram.vhd(68[19:45])
    defparam i1435_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2311_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_208_7), .O(n2559));   // src/ram.vhd(68[19:45])
    defparam i2311_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1434_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_99_2), .O(n1682));   // src/ram.vhd(68[19:45])
    defparam i1434_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1433_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_99_1), .O(n1681));   // src/ram.vhd(68[19:45])
    defparam i1433_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1587_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_118_3), .O(n1835));   // src/ram.vhd(68[19:45])
    defparam i1587_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2310_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_208_6), .O(n2558));   // src/ram.vhd(68[19:45])
    defparam i2310_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1432_3_lut_4_lut (.I0(n205), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_99_0), .O(n1680));   // src/ram.vhd(68[19:45])
    defparam i1432_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2391_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_218_7), .O(n2639));   // src/ram.vhd(68[19:45])
    defparam i2391_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2309_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_208_5), .O(n2557));   // src/ram.vhd(68[19:45])
    defparam i2309_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2390_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_218_6), .O(n2638));   // src/ram.vhd(68[19:45])
    defparam i2390_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2389_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_218_5), .O(n2637));   // src/ram.vhd(68[19:45])
    defparam i2389_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2388_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_218_4), .O(n2636));   // src/ram.vhd(68[19:45])
    defparam i2388_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2387_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_218_3), .O(n2635));   // src/ram.vhd(68[19:45])
    defparam i2387_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2386_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_218_2), .O(n2634));   // src/ram.vhd(68[19:45])
    defparam i2386_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1255_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_76_7), .O(n1503));   // src/ram.vhd(68[19:45])
    defparam i1255_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2308_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_208_4), .O(n2556));   // src/ram.vhd(68[19:45])
    defparam i2308_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2385_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_218_1), .O(n2633));   // src/ram.vhd(68[19:45])
    defparam i2385_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2384_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_218_0), .O(n2632));   // src/ram.vhd(68[19:45])
    defparam i2384_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2307_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_208_3), .O(n2555));   // src/ram.vhd(68[19:45])
    defparam i2307_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9204_3_lut (.I0(ram_s_152_7), .I1(ram_s_153_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10263));
    defparam i9204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9205_3_lut (.I0(ram_s_154_7), .I1(ram_s_155_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10264));
    defparam i9205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2306_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_208_2), .O(n2554));   // src/ram.vhd(68[19:45])
    defparam i2306_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9220_3_lut (.I0(ram_s_158_7), .I1(ram_s_159_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10279));
    defparam i9220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9219_3_lut (.I0(ram_s_156_7), .I1(ram_s_157_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10278));
    defparam i9219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8895_3_lut (.I0(ram_s_192_4), .I1(ram_s_193_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9954));
    defparam i8895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8896_3_lut (.I0(ram_s_194_4), .I1(ram_s_195_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9955));
    defparam i8896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1586_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_118_2), .O(n1834));   // src/ram.vhd(68[19:45])
    defparam i1586_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8908_3_lut (.I0(ram_s_198_4), .I1(ram_s_199_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9967));
    defparam i8908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8907_3_lut (.I0(ram_s_196_4), .I1(ram_s_197_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9966));
    defparam i8907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8202_3_lut (.I0(ram_s_224_0), .I1(ram_s_225_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9261));
    defparam i8202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8203_3_lut (.I0(ram_s_226_0), .I1(ram_s_227_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9262));
    defparam i8203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8224_3_lut (.I0(ram_s_230_0), .I1(ram_s_231_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9283));
    defparam i8224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8223_3_lut (.I0(ram_s_228_0), .I1(ram_s_229_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9282));
    defparam i8223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8244_3_lut (.I0(ram_s_240_0), .I1(ram_s_241_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9303));
    defparam i8244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1585_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_118_1), .O(n1833));   // src/ram.vhd(68[19:45])
    defparam i1585_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8245_3_lut (.I0(ram_s_242_0), .I1(ram_s_243_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9304));
    defparam i8245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8254_3_lut (.I0(ram_s_246_0), .I1(ram_s_247_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9313));
    defparam i8254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8253_3_lut (.I0(ram_s_244_0), .I1(ram_s_245_0), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9312));
    defparam i8253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1584_3_lut_4_lut (.I0(n243_adj_881), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_118_0), .O(n1832));   // src/ram.vhd(68[19:45])
    defparam i1584_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2305_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_208_1), .O(n2553));   // src/ram.vhd(68[19:45])
    defparam i2305_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i234_2_lut_3_lut (.I0(n41), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n234));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i234_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1431_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_98_7), .O(n1679));   // src/ram.vhd(68[19:45])
    defparam i1431_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i233_2_lut_3_lut (.I0(n41), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n233));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i233_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2567_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_240_7), .O(n2815));   // src/ram.vhd(68[19:45])
    defparam i2567_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1430_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_98_6), .O(n1678));   // src/ram.vhd(68[19:45])
    defparam i1430_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1254_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_76_6), .O(n1502));   // src/ram.vhd(68[19:45])
    defparam i1254_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2304_3_lut_4_lut (.I0(n167), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_208_0), .O(n2552));   // src/ram.vhd(68[19:45])
    defparam i2304_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2566_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_240_6), .O(n2814));   // src/ram.vhd(68[19:45])
    defparam i2566_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1429_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_98_5), .O(n1677));   // src/ram.vhd(68[19:45])
    defparam i1429_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2565_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_240_5), .O(n2813));   // src/ram.vhd(68[19:45])
    defparam i2565_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1279_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_79_7), .O(n1527));   // src/ram.vhd(68[19:45])
    defparam i1279_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1278_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_79_6), .O(n1526));   // src/ram.vhd(68[19:45])
    defparam i1278_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2564_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_240_4), .O(n2812));   // src/ram.vhd(68[19:45])
    defparam i2564_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1428_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_98_4), .O(n1676));   // src/ram.vhd(68[19:45])
    defparam i1428_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1427_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_98_3), .O(n1675));   // src/ram.vhd(68[19:45])
    defparam i1427_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1277_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_79_5), .O(n1525));   // src/ram.vhd(68[19:45])
    defparam i1277_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1253_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_76_5), .O(n1501));   // src/ram.vhd(68[19:45])
    defparam i1253_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2563_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_240_3), .O(n2811));   // src/ram.vhd(68[19:45])
    defparam i2563_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1426_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_98_2), .O(n1674));   // src/ram.vhd(68[19:45])
    defparam i1426_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i20_2_lut (.I0(n11), .I1(port_id[2]), .I2(wea[0]), 
            .I3(wea[0]), .O(n20));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i20_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1425_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_98_1), .O(n1673));   // src/ram.vhd(68[19:45])
    defparam i1425_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1424_3_lut_4_lut (.I0(n203), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_98_0), .O(n1672));   // src/ram.vhd(68[19:45])
    defparam i1424_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1423_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_97_7), .O(n1671));   // src/ram.vhd(68[19:45])
    defparam i1423_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i156_2_lut (.I0(n92_c), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n156));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i156_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1422_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_97_6), .O(n1670));   // src/ram.vhd(68[19:45])
    defparam i1422_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1421_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_97_5), .O(n1669));   // src/ram.vhd(68[19:45])
    defparam i1421_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1420_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_97_4), .O(n1668));   // src/ram.vhd(68[19:45])
    defparam i1420_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2562_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_240_2), .O(n2810));   // src/ram.vhd(68[19:45])
    defparam i2562_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2561_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_240_1), .O(n2809));   // src/ram.vhd(68[19:45])
    defparam i2561_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2560_3_lut_4_lut (.I0(n231), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_240_0), .O(n2808));   // src/ram.vhd(68[19:45])
    defparam i2560_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1583_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_117_7), .O(n1831));   // src/ram.vhd(68[19:45])
    defparam i1583_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1582_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_117_6), .O(n1830));   // src/ram.vhd(68[19:45])
    defparam i1582_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1581_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_117_5), .O(n1829));   // src/ram.vhd(68[19:45])
    defparam i1581_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1580_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_117_4), .O(n1828));   // src/ram.vhd(68[19:45])
    defparam i1580_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1579_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_117_3), .O(n1827));   // src/ram.vhd(68[19:45])
    defparam i1579_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1276_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_79_4), .O(n1524));   // src/ram.vhd(68[19:45])
    defparam i1276_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1275_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_79_3), .O(n1523));   // src/ram.vhd(68[19:45])
    defparam i1275_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1419_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_97_3), .O(n1667));   // src/ram.vhd(68[19:45])
    defparam i1419_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i377_378 (.Q(ram_s_15_1), .C(CLK_3P3_MHZ_c), .D(n913));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1578_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_117_2), .O(n1826));   // src/ram.vhd(68[19:45])
    defparam i1578_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1418_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_97_2), .O(n1666));   // src/ram.vhd(68[19:45])
    defparam i1418_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1577_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_117_1), .O(n1825));   // src/ram.vhd(68[19:45])
    defparam i1577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1274_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_79_2), .O(n1522));   // src/ram.vhd(68[19:45])
    defparam i1274_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1417_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_97_1), .O(n1665));   // src/ram.vhd(68[19:45])
    defparam i1417_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1576_3_lut_4_lut (.I0(n241), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_117_0), .O(n1824));   // src/ram.vhd(68[19:45])
    defparam i1576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1273_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_79_1), .O(n1521));   // src/ram.vhd(68[19:45])
    defparam i1273_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1416_3_lut_4_lut (.I0(n201), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_97_0), .O(n1664));   // src/ram.vhd(68[19:45])
    defparam i1416_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i232_2_lut_3_lut (.I0(n39), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n232));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i232_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1272_3_lut_4_lut (.I0(n165), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_79_0), .O(n1520));   // src/ram.vhd(68[19:45])
    defparam i1272_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2383_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_217_7), .O(n2631));   // src/ram.vhd(68[19:45])
    defparam i2383_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i231_2_lut_3_lut (.I0(n39), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n231));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i231_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i168_2_lut_3_lut (.I0(n39), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n168));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i168_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i2382_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_217_6), .O(n2630));   // src/ram.vhd(68[19:45])
    defparam i2382_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i167_2_lut_3_lut (.I0(n39), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n167));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i167_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2381_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_217_5), .O(n2629));   // src/ram.vhd(68[19:45])
    defparam i2381_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut (.I0(n16), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(wea[0]), .O(n39));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i39_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1271_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_78_7), .O(n1519));   // src/ram.vhd(68[19:45])
    defparam i1271_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2380_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_217_4), .O(n2628));   // src/ram.vhd(68[19:45])
    defparam i2380_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i71_2_lut_3_lut_4_lut (.I0(n16), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n71_adj_842));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i71_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1270_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_78_6), .O(n1518));   // src/ram.vhd(68[19:45])
    defparam i1270_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2379_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_217_3), .O(n2627));   // src/ram.vhd(68[19:45])
    defparam i2379_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i72_2_lut_3_lut_4_lut (.I0(n16), .I1(port_id[3]), 
            .I2(port_id[5]), .I3(port_id[4]), .O(n72_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i72_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1269_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_78_5), .O(n1517));   // src/ram.vhd(68[19:45])
    defparam i1269_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2378_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_217_2), .O(n2626));   // src/ram.vhd(68[19:45])
    defparam i2378_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2559_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_239_7), .O(n2807));   // src/ram.vhd(68[19:45])
    defparam i2559_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1268_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_78_4), .O(n1516));   // src/ram.vhd(68[19:45])
    defparam i1268_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8268_3_lut (.I0(ram_s_72_6), .I1(ram_s_73_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9327));
    defparam i8268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8269_3_lut (.I0(ram_s_74_6), .I1(ram_s_75_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9328));
    defparam i8269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2377_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_217_1), .O(n2625));   // src/ram.vhd(68[19:45])
    defparam i2377_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1252_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_76_4), .O(n1500));   // src/ram.vhd(68[19:45])
    defparam i1252_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2558_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_239_6), .O(n2806));   // src/ram.vhd(68[19:45])
    defparam i2558_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11478 (.I0(port_id[0]), .I1(ram_s_254_4), 
            .I2(ram_s_255_4), .I3(port_id[1]), .O(n12809));
    defparam port_id_0__bdd_4_lut_11478.LUT_INIT = 16'he4aa;
    SB_LUT4 n12809_bdd_4_lut (.I0(n12809), .I1(ram_s_253_4), .I2(ram_s_252_4), 
            .I3(port_id[1]), .O(n12812));
    defparam n12809_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11518 (.I0(port_id[2]), .I1(n10640), .I2(n10664), 
            .I3(port_id[3]), .O(n12803));
    defparam port_id_2__bdd_4_lut_11518.LUT_INIT = 16'he4aa;
    SB_LUT4 n12803_bdd_4_lut (.I0(n12803), .I1(n10595), .I2(n10574), .I3(port_id[3]), 
            .O(n12806));
    defparam n12803_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11468 (.I0(port_id[0]), .I1(ram_s_118_2), 
            .I2(ram_s_119_2), .I3(port_id[1]), .O(n12797));
    defparam port_id_0__bdd_4_lut_11468.LUT_INIT = 16'he4aa;
    SB_LUT4 n12797_bdd_4_lut (.I0(n12797), .I1(ram_s_117_2), .I2(ram_s_116_2), 
            .I3(port_id[1]), .O(n12800));
    defparam n12797_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2376_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_217_0), .O(n2624));   // src/ram.vhd(68[19:45])
    defparam i2376_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11458 (.I0(port_id[0]), .I1(ram_s_82_4), 
            .I2(ram_s_83_4), .I3(port_id[1]), .O(n12791));
    defparam port_id_0__bdd_4_lut_11458.LUT_INIT = 16'he4aa;
    SB_LUT4 n12791_bdd_4_lut (.I0(n12791), .I1(ram_s_81_4), .I2(ram_s_80_4), 
            .I3(port_id[1]), .O(n9710));
    defparam n12791_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11453 (.I0(port_id[0]), .I1(ram_s_10_5), 
            .I2(ram_s_11_5), .I3(port_id[1]), .O(n12785));
    defparam port_id_0__bdd_4_lut_11453.LUT_INIT = 16'he4aa;
    SB_LUT4 n12785_bdd_4_lut (.I0(n12785), .I1(ram_s_9_5), .I2(ram_s_8_5), 
            .I3(port_id[1]), .O(n10826));
    defparam n12785_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11448 (.I0(port_id[0]), .I1(ram_s_78_7), 
            .I2(ram_s_79_7), .I3(port_id[1]), .O(n12773));
    defparam port_id_0__bdd_4_lut_11448.LUT_INIT = 16'he4aa;
    SB_LUT4 n12773_bdd_4_lut (.I0(n12773), .I1(ram_s_77_7), .I2(ram_s_76_7), 
            .I3(port_id[1]), .O(n12776));
    defparam n12773_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11438 (.I0(port_id[0]), .I1(ram_s_106_3), 
            .I2(ram_s_107_3), .I3(port_id[1]), .O(n12767));
    defparam port_id_0__bdd_4_lut_11438.LUT_INIT = 16'he4aa;
    SB_LUT4 n12767_bdd_4_lut (.I0(n12767), .I1(ram_s_105_3), .I2(ram_s_104_3), 
            .I3(port_id[1]), .O(n9368));
    defparam n12767_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11433 (.I0(port_id[0]), .I1(ram_s_18_6), 
            .I2(ram_s_19_6), .I3(port_id[1]), .O(n12761));
    defparam port_id_0__bdd_4_lut_11433.LUT_INIT = 16'he4aa;
    SB_LUT4 n12761_bdd_4_lut (.I0(n12761), .I1(ram_s_17_6), .I2(ram_s_16_6), 
            .I3(port_id[1]), .O(n9074));
    defparam n12761_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2557_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_239_5), .O(n2805));   // src/ram.vhd(68[19:45])
    defparam i2557_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2556_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_239_4), .O(n2804));   // src/ram.vhd(68[19:45])
    defparam i2556_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2555_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_239_3), .O(n2803));   // src/ram.vhd(68[19:45])
    defparam i2555_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11428 (.I0(port_id[0]), .I1(ram_s_142_1), 
            .I2(ram_s_143_1), .I3(port_id[1]), .O(n12755));
    defparam port_id_0__bdd_4_lut_11428.LUT_INIT = 16'he4aa;
    SB_LUT4 i8278_3_lut (.I0(ram_s_78_6), .I1(ram_s_79_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9337));
    defparam i8278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12755_bdd_4_lut (.I0(n12755), .I1(ram_s_141_1), .I2(ram_s_140_1), 
            .I3(port_id[1]), .O(n12758));
    defparam n12755_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11423 (.I0(port_id[0]), .I1(ram_s_6_1), 
            .I2(ram_s_7_1), .I3(port_id[1]), .O(n12749));
    defparam port_id_0__bdd_4_lut_11423.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11050 (.I0(port_id[0]), .I1(ram_s_22_1), 
            .I2(ram_s_23_1), .I3(port_id[1]), .O(n12299));
    defparam port_id_0__bdd_4_lut_11050.LUT_INIT = 16'he4aa;
    SB_LUT4 n12749_bdd_4_lut (.I0(n12749), .I1(ram_s_5_1), .I2(ram_s_4_1), 
            .I3(port_id[1]), .O(n12752));
    defparam n12749_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12299_bdd_4_lut (.I0(n12299), .I1(ram_s_21_1), .I2(ram_s_20_1), 
            .I3(port_id[1]), .O(n12302));
    defparam n12299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8277_3_lut (.I0(ram_s_76_6), .I1(ram_s_77_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9336));
    defparam i8277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2375_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_216_7), .O(n2623));   // src/ram.vhd(68[19:45])
    defparam i2375_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_2__bdd_4_lut_11463 (.I0(port_id[2]), .I1(n10676), .I2(n10679), 
            .I3(port_id[3]), .O(n12743));
    defparam port_id_2__bdd_4_lut_11463.LUT_INIT = 16'he4aa;
    SB_LUT4 n12743_bdd_4_lut (.I0(n12743), .I1(n10667), .I2(n10658), .I3(port_id[3]), 
            .O(n10829));
    defparam n12743_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11418 (.I0(port_id[0]), .I1(ram_s_74_5), 
            .I2(ram_s_75_5), .I3(port_id[1]), .O(n12737));
    defparam port_id_0__bdd_4_lut_11418.LUT_INIT = 16'he4aa;
    SB_LUT4 n12737_bdd_4_lut (.I0(n12737), .I1(ram_s_73_5), .I2(ram_s_72_5), 
            .I3(port_id[1]), .O(n12740));
    defparam n12737_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11408 (.I0(port_id[0]), .I1(ram_s_86_4), 
            .I2(ram_s_87_4), .I3(port_id[1]), .O(n12731));
    defparam port_id_0__bdd_4_lut_11408.LUT_INIT = 16'he4aa;
    SB_LUT4 n12731_bdd_4_lut (.I0(n12731), .I1(ram_s_85_4), .I2(ram_s_84_4), 
            .I3(port_id[1]), .O(n9719));
    defparam n12731_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11045 (.I0(port_id[0]), .I1(ram_s_254_5), 
            .I2(ram_s_255_5), .I3(port_id[1]), .O(n12293));
    defparam port_id_0__bdd_4_lut_11045.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10890 (.I0(port_id[2]), .I1(n10412), .I2(n10427), 
            .I3(port_id[3]), .O(n12077));
    defparam port_id_2__bdd_4_lut_10890.LUT_INIT = 16'he4aa;
    SB_LUT4 i1251_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_76_3), .O(n1499));   // src/ram.vhd(68[19:45])
    defparam i1251_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12077_bdd_4_lut (.I0(n12077), .I1(n10394), .I2(n10370), .I3(port_id[3]), 
            .O(n12080));
    defparam n12077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11693_bdd_4_lut (.I0(n11693), .I1(ram_s_189_1), .I2(ram_s_188_1), 
            .I3(port_id[1]), .O(n11696));
    defparam n11693_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10700 (.I0(port_id[2]), .I1(n9119), .I2(n9131), 
            .I3(port_id[3]), .O(n11873));
    defparam port_id_2__bdd_4_lut_10700.LUT_INIT = 16'he4aa;
    SB_LUT4 i2554_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_239_2), .O(n2802));   // src/ram.vhd(68[19:45])
    defparam i2554_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2374_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_216_6), .O(n2622));   // src/ram.vhd(68[19:45])
    defparam i2374_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2553_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_239_1), .O(n2801));   // src/ram.vhd(68[19:45])
    defparam i2553_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11873_bdd_4_lut (.I0(n11873), .I1(n9101), .I2(n9074), .I3(port_id[3]), 
            .O(n11876));
    defparam n11873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10431 (.I0(port_id[0]), .I1(ram_s_182_6), 
            .I2(ram_s_183_6), .I3(port_id[1]), .O(n11543));
    defparam port_id_0__bdd_4_lut_10431.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10860 (.I0(port_id[2]), .I1(n9227), .I2(n9251), 
            .I3(port_id[3]), .O(n12071));
    defparam port_id_2__bdd_4_lut_10860.LUT_INIT = 16'he4aa;
    SB_LUT4 i2373_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_216_5), .O(n2621));   // src/ram.vhd(68[19:45])
    defparam i2373_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12071_bdd_4_lut (.I0(n12071), .I1(n9182), .I2(n9161), .I3(port_id[3]), 
            .O(n12074));
    defparam n12071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12293_bdd_4_lut (.I0(n12293), .I1(ram_s_253_5), .I2(ram_s_252_5), 
            .I3(port_id[1]), .O(n10475));
    defparam n12293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11543_bdd_4_lut (.I0(n11543), .I1(ram_s_181_6), .I2(ram_s_180_6), 
            .I3(port_id[1]), .O(n11546));
    defparam n11543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2372_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_216_4), .O(n2620));   // src/ram.vhd(68[19:45])
    defparam i2372_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_4__bdd_4_lut_11025 (.I0(port_id[4]), .I1(n11009), .I2(n11015), 
            .I3(port_id[5]), .O(n11687));
    defparam port_id_4__bdd_4_lut_11025.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10745 (.I0(port_id[0]), .I1(ram_s_254_6), 
            .I2(ram_s_255_6), .I3(port_id[1]), .O(n11867));
    defparam port_id_0__bdd_4_lut_10745.LUT_INIT = 16'he4aa;
    SB_LUT4 n11687_bdd_4_lut (.I0(n11687), .I1(n11540), .I2(n11060), .I3(port_id[5]), 
            .O(n11690));
    defparam n11687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11867_bdd_4_lut (.I0(n11867), .I1(ram_s_253_6), .I2(ram_s_252_6), 
            .I3(port_id[1]), .O(n11870));
    defparam n11867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10865 (.I0(port_id[0]), .I1(ram_s_22_0), 
            .I2(ram_s_23_0), .I3(port_id[1]), .O(n12065));
    defparam port_id_0__bdd_4_lut_10865.LUT_INIT = 16'he4aa;
    SB_LUT4 n12065_bdd_4_lut (.I0(n12065), .I1(ram_s_21_0), .I2(ram_s_20_0), 
            .I3(port_id[1]), .O(n12068));
    defparam n12065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10591 (.I0(port_id[2]), .I1(n9068), .I2(n9077), 
            .I3(port_id[3]), .O(n11681));
    defparam port_id_2__bdd_4_lut_10591.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10850 (.I0(port_id[0]), .I1(ram_s_114_5), 
            .I2(ram_s_115_5), .I3(port_id[1]), .O(n12059));
    defparam port_id_0__bdd_4_lut_10850.LUT_INIT = 16'he4aa;
    SB_LUT4 n11681_bdd_4_lut (.I0(n11681), .I1(n9065), .I2(n9053), .I3(port_id[3]), 
            .O(n11684));
    defparam n11681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2371_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_216_3), .O(n2619));   // src/ram.vhd(68[19:45])
    defparam i2371_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2370_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_216_2), .O(n2618));   // src/ram.vhd(68[19:45])
    defparam i2370_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_2__bdd_4_lut_10426 (.I0(port_id[2]), .I1(n9728), .I2(n9737), 
            .I3(port_id[3]), .O(n11537));
    defparam port_id_2__bdd_4_lut_10426.LUT_INIT = 16'he4aa;
    SB_LUT4 n12059_bdd_4_lut (.I0(n12059), .I1(ram_s_113_5), .I2(ram_s_112_5), 
            .I3(port_id[1]), .O(n12062));
    defparam n12059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8386_3_lut (.I0(n14450), .I1(n14348), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9445));
    defparam i8386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 port_id_0__bdd_4_lut_11040 (.I0(port_id[0]), .I1(ram_s_138_5), 
            .I2(ram_s_139_5), .I3(port_id[1]), .O(n12287));
    defparam port_id_0__bdd_4_lut_11040.LUT_INIT = 16'he4aa;
    SB_LUT4 n12287_bdd_4_lut (.I0(n12287), .I1(ram_s_137_5), .I2(ram_s_136_5), 
            .I3(port_id[1]), .O(n12290));
    defparam n12287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2369_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_216_1), .O(n2617));   // src/ram.vhd(68[19:45])
    defparam i2369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10845 (.I0(port_id[0]), .I1(ram_s_38_2), 
            .I2(ram_s_39_2), .I3(port_id[1]), .O(n12053));
    defparam port_id_0__bdd_4_lut_10845.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10690 (.I0(port_id[2]), .I1(n9905), .I2(n9917), 
            .I3(port_id[3]), .O(n11855));
    defparam port_id_2__bdd_4_lut_10690.LUT_INIT = 16'he4aa;
    SB_LUT4 n11855_bdd_4_lut (.I0(n11855), .I1(n9899), .I2(n9884), .I3(port_id[3]), 
            .O(n11054));
    defparam n11855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11403 (.I0(port_id[0]), .I1(ram_s_146_1), 
            .I2(ram_s_147_1), .I3(port_id[1]), .O(n12719));
    defparam port_id_0__bdd_4_lut_11403.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_1__bdd_4_lut_10950 (.I0(port_id[1]), .I1(n10065), .I2(n10066), 
            .I3(port_id[2]), .O(n11849));
    defparam port_id_1__bdd_4_lut_10950.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11035 (.I0(port_id[0]), .I1(ram_s_198_3), 
            .I2(ram_s_199_3), .I3(port_id[1]), .O(n12281));
    defparam port_id_0__bdd_4_lut_11035.LUT_INIT = 16'he4aa;
    SB_LUT4 n12053_bdd_4_lut (.I0(n12053), .I1(ram_s_37_2), .I2(ram_s_36_2), 
            .I3(port_id[1]), .O(n12056));
    defparam n12053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12281_bdd_4_lut (.I0(n12281), .I1(ram_s_197_3), .I2(ram_s_196_3), 
            .I3(port_id[1]), .O(n12284));
    defparam n12281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11849_bdd_4_lut (.I0(n11849), .I1(n10048), .I2(n10047), .I3(port_id[2]), 
            .O(n11852));
    defparam n11849_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10541 (.I0(port_id[0]), .I1(ram_s_74_3), 
            .I2(ram_s_75_3), .I3(port_id[1]), .O(n11675));
    defparam port_id_0__bdd_4_lut_10541.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_4__bdd_4_lut_11169 (.I0(port_id[4]), .I1(n9278), .I2(n9941), 
            .I3(port_id[5]), .O(n12275));
    defparam port_id_4__bdd_4_lut_11169.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10840 (.I0(port_id[0]), .I1(ram_s_46_5), 
            .I2(ram_s_47_5), .I3(port_id[1]), .O(n12047));
    defparam port_id_0__bdd_4_lut_10840.LUT_INIT = 16'he4aa;
    SB_LUT4 n12047_bdd_4_lut (.I0(n12047), .I1(ram_s_45_5), .I2(ram_s_44_5), 
            .I3(port_id[1]), .O(n12050));
    defparam n12047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12275_bdd_4_lut (.I0(n12275), .I1(n8825), .I2(n10646), .I3(port_id[5]), 
            .O(n12278));
    defparam n12275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11030 (.I0(port_id[0]), .I1(ram_s_6_0), 
            .I2(ram_s_7_0), .I3(port_id[1]), .O(n12269));
    defparam port_id_0__bdd_4_lut_11030.LUT_INIT = 16'he4aa;
    SB_LUT4 n12269_bdd_4_lut (.I0(n12269), .I1(ram_s_5_0), .I2(ram_s_4_0), 
            .I3(port_id[1]), .O(n12272));
    defparam n12269_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11675_bdd_4_lut (.I0(n11675), .I1(ram_s_73_3), .I2(ram_s_72_3), 
            .I3(port_id[1]), .O(n11678));
    defparam n11675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11020 (.I0(port_id[0]), .I1(ram_s_162_1), 
            .I2(ram_s_163_1), .I3(port_id[1]), .O(n12263));
    defparam port_id_0__bdd_4_lut_11020.LUT_INIT = 16'he4aa;
    SB_LUT4 n11537_bdd_4_lut (.I0(n11537), .I1(n9719), .I2(n9710), .I3(port_id[3]), 
            .O(n11540));
    defparam n11537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12719_bdd_4_lut (.I0(n12719), .I1(ram_s_145_1), .I2(ram_s_144_1), 
            .I3(port_id[1]), .O(n12722));
    defparam n12719_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11393 (.I0(port_id[0]), .I1(ram_s_190_3), 
            .I2(ram_s_191_3), .I3(port_id[1]), .O(n12713));
    defparam port_id_0__bdd_4_lut_11393.LUT_INIT = 16'he4aa;
    SB_LUT4 n12713_bdd_4_lut (.I0(n12713), .I1(ram_s_189_3), .I2(ram_s_188_3), 
            .I3(port_id[1]), .O(n12716));
    defparam n12713_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2368_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_216_0), .O(n2616));   // src/ram.vhd(68[19:45])
    defparam i2368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11388 (.I0(port_id[0]), .I1(ram_s_142_0), 
            .I2(ram_s_143_0), .I3(port_id[1]), .O(n12707));
    defparam port_id_0__bdd_4_lut_11388.LUT_INIT = 16'he4aa;
    SB_LUT4 n12707_bdd_4_lut (.I0(n12707), .I1(ram_s_141_0), .I2(ram_s_140_0), 
            .I3(port_id[1]), .O(n9077));
    defparam n12707_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11538 (.I0(port_id[1]), .I1(n9564), .I2(n9565), 
            .I3(port_id[2]), .O(n12701));
    defparam port_id_1__bdd_4_lut_11538.LUT_INIT = 16'he4aa;
    SB_LUT4 n12701_bdd_4_lut (.I0(n12701), .I1(n9547), .I2(n9546), .I3(port_id[2]), 
            .O(n10102));
    defparam n12701_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11383 (.I0(port_id[0]), .I1(ram_s_14_2), 
            .I2(ram_s_15_2), .I3(port_id[1]), .O(n12695));
    defparam port_id_0__bdd_4_lut_11383.LUT_INIT = 16'he4aa;
    SB_LUT4 n12695_bdd_4_lut (.I0(n12695), .I1(ram_s_13_2), .I2(ram_s_12_2), 
            .I3(port_id[1]), .O(n12698));
    defparam n12695_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11413 (.I0(port_id[2]), .I1(n12380), .I2(n12242), 
            .I3(port_id[3]), .O(n12689));
    defparam port_id_2__bdd_4_lut_11413.LUT_INIT = 16'he4aa;
    SB_LUT4 n12689_bdd_4_lut (.I0(n12689), .I1(n12440), .I2(n12626), .I3(port_id[3]), 
            .O(n12692));
    defparam n12689_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12263_bdd_4_lut (.I0(n12263), .I1(ram_s_161_1), .I2(ram_s_160_1), 
            .I3(port_id[1]), .O(n12266));
    defparam n12263_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10835 (.I0(port_id[0]), .I1(ram_s_46_3), 
            .I2(ram_s_47_3), .I3(port_id[1]), .O(n12041));
    defparam port_id_0__bdd_4_lut_10835.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10526 (.I0(port_id[0]), .I1(ram_s_194_5), 
            .I2(ram_s_195_5), .I3(port_id[1]), .O(n11669));
    defparam port_id_0__bdd_4_lut_10526.LUT_INIT = 16'he4aa;
    SB_LUT4 i1267_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_78_3), .O(n1515));   // src/ram.vhd(68[19:45])
    defparam i1267_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i184_2_lut_3_lut (.I0(n55_adj_879), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n184_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i184_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1266_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_78_2), .O(n1514));   // src/ram.vhd(68[19:45])
    defparam i1266_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2552_3_lut_4_lut (.I0(n229), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_239_0), .O(n2800));   // src/ram.vhd(68[19:45])
    defparam i2552_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11669_bdd_4_lut (.I0(n11669), .I1(ram_s_193_5), .I2(ram_s_192_5), 
            .I3(port_id[1]), .O(n11672));
    defparam n11669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i521_522 (.Q(ram_s_21_1), .C(CLK_3P3_MHZ_c), .D(n912));   // src/ram.vhd(56[12:17])
    SB_LUT4 i8392_3_lut (.I0(n14090), .I1(n14006), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9451));
    defparam i8392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i183_2_lut_3_lut (.I0(n55_adj_879), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n183_adj_883));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i183_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1265_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_78_1), .O(n1513));   // src/ram.vhd(68[19:45])
    defparam i1265_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1415_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_96_7), .O(n1663));   // src/ram.vhd(68[19:45])
    defparam i1415_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1414_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_96_6), .O(n1662));   // src/ram.vhd(68[19:45])
    defparam i1414_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12041_bdd_4_lut (.I0(n12041), .I1(ram_s_45_3), .I2(ram_s_44_3), 
            .I3(port_id[1]), .O(n12044));
    defparam n12041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11368 (.I0(port_id[2]), .I1(n9959), .I2(n9980), 
            .I3(port_id[3]), .O(n12677));
    defparam port_id_2__bdd_4_lut_11368.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i165_2_lut_3_lut_4_lut (.I0(n37), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n165));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i165_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i8424_3_lut (.I0(n13124), .I1(n13016), .I2(port_id[4]), .I3(wea[0]), 
            .O(n9483));
    defparam i8424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1413_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_96_5), .O(n1661));   // src/ram.vhd(68[19:45])
    defparam i1413_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_2__bdd_4_lut_10675 (.I0(port_id[2]), .I1(n9692), .I2(n9707), 
            .I3(port_id[3]), .O(n11837));
    defparam port_id_2__bdd_4_lut_10675.LUT_INIT = 16'he4aa;
    SB_LUT4 i8425_3_lut (.I0(n12884), .I1(n12872), .I2(port_id[4]), .I3(wea[0]), 
            .O(n9484));
    defparam i8425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 port_id_2__bdd_4_lut_10531 (.I0(port_id[2]), .I1(n9512), .I2(n9536), 
            .I3(port_id[3]), .O(n11663));
    defparam port_id_2__bdd_4_lut_10531.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i166_2_lut_3_lut_4_lut (.I0(n37), .I1(port_id[4]), 
            .I2(port_id[6]), .I3(port_id[5]), .O(n166));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i166_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 port_id_0__bdd_4_lut_10830 (.I0(port_id[0]), .I1(ram_s_178_1), 
            .I2(ram_s_179_1), .I3(port_id[1]), .O(n12035));
    defparam port_id_0__bdd_4_lut_10830.LUT_INIT = 16'he4aa;
    SB_LUT4 n11837_bdd_4_lut (.I0(n11837), .I1(n9686), .I2(n9674), .I3(port_id[3]), 
            .O(n11060));
    defparam n11837_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10417 (.I0(port_id[0]), .I1(ram_s_118_5), 
            .I2(ram_s_119_5), .I3(port_id[1]), .O(n11531));
    defparam port_id_0__bdd_4_lut_10417.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11015 (.I0(port_id[0]), .I1(ram_s_10_0), 
            .I2(ram_s_11_0), .I3(port_id[1]), .O(n12257));
    defparam port_id_0__bdd_4_lut_11015.LUT_INIT = 16'he4aa;
    SB_LUT4 n11663_bdd_4_lut (.I0(n11663), .I1(n9461), .I2(n9440), .I3(port_id[3]), 
            .O(n11666));
    defparam n11663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1575_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_116_7), .O(n1823));   // src/ram.vhd(68[19:45])
    defparam i1575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12035_bdd_4_lut (.I0(n12035), .I1(ram_s_177_1), .I2(ram_s_176_1), 
            .I3(port_id[1]), .O(n12038));
    defparam n12035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1574_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_116_6), .O(n1822));   // src/ram.vhd(68[19:45])
    defparam i1574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12677_bdd_4_lut (.I0(n12677), .I1(n9923), .I2(n9887), .I3(port_id[3]), 
            .O(n12680));
    defparam n12677_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8437_3_lut (.I0(n12218), .I1(n12014), .I2(port_id[4]), .I3(wea[0]), 
            .O(n9496));
    defparam i8437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8436_3_lut (.I0(n12674), .I1(n12578), .I2(port_id[4]), .I3(wea[0]), 
            .O(n9495));
    defparam i8436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1412_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_96_4), .O(n1660));   // src/ram.vhd(68[19:45])
    defparam i1412_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1573_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_116_5), .O(n1821));   // src/ram.vhd(68[19:45])
    defparam i1573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1572_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_116_4), .O(n1820));   // src/ram.vhd(68[19:45])
    defparam i1572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1571_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_116_3), .O(n1819));   // src/ram.vhd(68[19:45])
    defparam i1571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_2__bdd_4_lut_11358 (.I0(port_id[2]), .I1(n8930), .I2(n8939), 
            .I3(port_id[3]), .O(n12671));
    defparam port_id_2__bdd_4_lut_11358.LUT_INIT = 16'he4aa;
    SB_LUT4 n12671_bdd_4_lut (.I0(n12671), .I1(n8927), .I2(n11510), .I3(port_id[3]), 
            .O(n12674));
    defparam n12671_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1411_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_96_3), .O(n1659));   // src/ram.vhd(68[19:45])
    defparam i1411_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1410_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_96_2), .O(n1658));   // src/ram.vhd(68[19:45])
    defparam i1410_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1570_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_116_2), .O(n1818));   // src/ram.vhd(68[19:45])
    defparam i1570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11373 (.I0(port_id[0]), .I1(ram_s_146_3), 
            .I2(ram_s_147_3), .I3(port_id[1]), .O(n12665));
    defparam port_id_0__bdd_4_lut_11373.LUT_INIT = 16'he4aa;
    SB_LUT4 n12665_bdd_4_lut (.I0(n12665), .I1(ram_s_145_3), .I2(ram_s_144_3), 
            .I3(port_id[1]), .O(n9725));
    defparam n12665_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1264_3_lut_4_lut (.I0(n163), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_78_0), .O(n1512));   // src/ram.vhd(68[19:45])
    defparam i1264_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1569_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_116_1), .O(n1817));   // src/ram.vhd(68[19:45])
    defparam i1569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1409_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_96_1), .O(n1657));   // src/ram.vhd(68[19:45])
    defparam i1409_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1568_3_lut_4_lut (.I0(n239), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_116_0), .O(n1816));   // src/ram.vhd(68[19:45])
    defparam i1568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_11348 (.I0(port_id[0]), .I1(ram_s_90_4), 
            .I2(ram_s_91_4), .I3(port_id[1]), .O(n12659));
    defparam port_id_0__bdd_4_lut_11348.LUT_INIT = 16'he4aa;
    SB_DFF i332_333 (.Q(ram_s_13_2), .C(CLK_3P3_MHZ_c), .D(n911));   // src/ram.vhd(56[12:17])
    SB_DFF i275_276 (.Q(ram_s_10_7), .C(CLK_3P3_MHZ_c), .D(n910));   // src/ram.vhd(56[12:17])
    SB_DFF i278_279 (.Q(ram_s_11_0), .C(CLK_3P3_MHZ_c), .D(n909));   // src/ram.vhd(56[12:17])
    SB_DFF i359_360 (.Q(ram_s_14_3), .C(CLK_3P3_MHZ_c), .D(n908));   // src/ram.vhd(56[12:17])
    SB_DFF i329_330 (.Q(ram_s_13_1), .C(CLK_3P3_MHZ_c), .D(n907));   // src/ram.vhd(56[12:17])
    SB_DFF i356_357 (.Q(ram_s_14_2), .C(CLK_3P3_MHZ_c), .D(n906));   // src/ram.vhd(56[12:17])
    SB_LUT4 i1408_3_lut_4_lut (.I0(n199_adj_843), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_96_0), .O(n1656));   // src/ram.vhd(68[19:45])
    defparam i1408_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i524_525 (.Q(ram_s_21_2), .C(CLK_3P3_MHZ_c), .D(n905));   // src/ram.vhd(56[12:17])
    SB_DFF i326_327 (.Q(ram_s_13_0), .C(CLK_3P3_MHZ_c), .D(n904));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2551_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_238_7), .O(n2799));   // src/ram.vhd(68[19:45])
    defparam i2551_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i380_381 (.Q(ram_s_15_2), .C(CLK_3P3_MHZ_c), .D(n903));   // src/ram.vhd(56[12:17])
    SB_DFF i383_384 (.Q(ram_s_15_3), .C(CLK_3P3_MHZ_c), .D(n902));   // src/ram.vhd(56[12:17])
    SB_DFF i146_147 (.Q(ram_s_5_4), .C(CLK_3P3_MHZ_c), .D(n901));   // src/ram.vhd(56[12:17])
    SB_DFF i386_387 (.Q(ram_s_15_4), .C(CLK_3P3_MHZ_c), .D(n900));   // src/ram.vhd(56[12:17])
    SB_DFF i368_369 (.Q(ram_s_14_6), .C(CLK_3P3_MHZ_c), .D(n899));   // src/ram.vhd(56[12:17])
    SB_LUT4 i2550_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_238_6), .O(n2798));   // src/ram.vhd(68[19:45])
    defparam i2550_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12659_bdd_4_lut (.I0(n12659), .I1(ram_s_89_4), .I2(ram_s_88_4), 
            .I3(port_id[1]), .O(n9728));
    defparam n12659_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2549_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_238_5), .O(n2797));   // src/ram.vhd(68[19:45])
    defparam i2549_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1263_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_77_7), .O(n1511));   // src/ram.vhd(68[19:45])
    defparam i1263_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1407_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_95_7), .O(n1655));   // src/ram.vhd(68[19:45])
    defparam i1407_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1406_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_95_6), .O(n1654));   // src/ram.vhd(68[19:45])
    defparam i1406_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1405_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_95_5), .O(n1653));   // src/ram.vhd(68[19:45])
    defparam i1405_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_1__bdd_4_lut_11378 (.I0(port_id[1]), .I1(n9594), .I2(n9595), 
            .I3(port_id[2]), .O(n12653));
    defparam port_id_1__bdd_4_lut_11378.LUT_INIT = 16'he4aa;
    SB_LUT4 n12653_bdd_4_lut (.I0(n12653), .I1(n9586), .I2(n9585), .I3(port_id[2]), 
            .O(n10105));
    defparam n12653_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_11973 (.I0(port_id[4]), .I1(n10712), .I2(n10715), 
            .I3(port_id[5]), .O(n12647));
    defparam port_id_4__bdd_4_lut_11973.LUT_INIT = 16'he4aa;
    SB_LUT4 n12647_bdd_4_lut (.I0(n12647), .I1(n10703), .I2(n10694), .I3(port_id[5]), 
            .O(n10838));
    defparam n12647_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11343 (.I0(port_id[0]), .I1(ram_s_250_5), 
            .I2(ram_s_251_5), .I3(port_id[1]), .O(n12641));
    defparam port_id_0__bdd_4_lut_11343.LUT_INIT = 16'he4aa;
    SB_LUT4 n12641_bdd_4_lut (.I0(n12641), .I1(ram_s_249_5), .I2(ram_s_248_5), 
            .I3(port_id[1]), .O(n10439));
    defparam n12641_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11328 (.I0(port_id[0]), .I1(ram_s_170_6), 
            .I2(ram_s_171_6), .I3(port_id[1]), .O(n12635));
    defparam port_id_0__bdd_4_lut_11328.LUT_INIT = 16'he4aa;
    SB_LUT4 n12635_bdd_4_lut (.I0(n12635), .I1(ram_s_169_6), .I2(ram_s_168_6), 
            .I3(port_id[1]), .O(n12638));
    defparam n12635_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11353 (.I0(port_id[2]), .I1(n11750), .I2(n11480), 
            .I3(port_id[3]), .O(n12629));
    defparam port_id_2__bdd_4_lut_11353.LUT_INIT = 16'he4aa;
    SB_LUT4 n12629_bdd_4_lut (.I0(n12629), .I1(n12056), .I2(n12092), .I3(port_id[3]), 
            .O(n12632));
    defparam n12629_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10825 (.I0(port_id[0]), .I1(ram_s_26_0), 
            .I2(ram_s_27_0), .I3(port_id[1]), .O(n12029));
    defparam port_id_0__bdd_4_lut_10825.LUT_INIT = 16'he4aa;
    SB_LUT4 n12257_bdd_4_lut (.I0(n12257), .I1(ram_s_9_0), .I2(ram_s_8_0), 
            .I3(port_id[1]), .O(n12260));
    defparam n12257_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11531_bdd_4_lut (.I0(n11531), .I1(ram_s_117_5), .I2(ram_s_116_5), 
            .I3(port_id[1]), .O(n11534));
    defparam n11531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11323 (.I0(port_id[0]), .I1(ram_s_18_2), 
            .I2(ram_s_19_2), .I3(port_id[1]), .O(n12623));
    defparam port_id_0__bdd_4_lut_11323.LUT_INIT = 16'he4aa;
    SB_LUT4 n12623_bdd_4_lut (.I0(n12623), .I1(ram_s_17_2), .I2(ram_s_16_2), 
            .I3(port_id[1]), .O(n12626));
    defparam n12623_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12029_bdd_4_lut (.I0(n12029), .I1(ram_s_25_0), .I2(ram_s_24_0), 
            .I3(port_id[1]), .O(n12032));
    defparam n12029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10820 (.I0(port_id[0]), .I1(ram_s_210_7), 
            .I2(ram_s_211_7), .I3(port_id[1]), .O(n12023));
    defparam port_id_0__bdd_4_lut_10820.LUT_INIT = 16'he4aa;
    SB_LUT4 n12023_bdd_4_lut (.I0(n12023), .I1(ram_s_209_7), .I2(ram_s_208_7), 
            .I3(port_id[1]), .O(n10517));
    defparam n12023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11010 (.I0(port_id[0]), .I1(ram_s_202_7), 
            .I2(ram_s_203_7), .I3(port_id[1]), .O(n12251));
    defparam port_id_0__bdd_4_lut_11010.LUT_INIT = 16'he4aa;
    SB_LUT4 i1404_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_95_4), .O(n1652));   // src/ram.vhd(68[19:45])
    defparam i1404_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_2__bdd_4_lut_10660 (.I0(port_id[2]), .I1(n9944), .I2(n9953), 
            .I3(port_id[3]), .O(n11819));
    defparam port_id_2__bdd_4_lut_10660.LUT_INIT = 16'he4aa;
    SB_LUT4 n11819_bdd_4_lut (.I0(n11819), .I1(n9929), .I2(n9920), .I3(port_id[3]), 
            .O(n11072));
    defparam n11819_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12251_bdd_4_lut (.I0(n12251), .I1(ram_s_201_7), .I2(ram_s_200_7), 
            .I3(port_id[1]), .O(n10481));
    defparam n12251_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11313 (.I0(port_id[0]), .I1(ram_s_110_5), 
            .I2(ram_s_111_5), .I3(port_id[1]), .O(n12617));
    defparam port_id_0__bdd_4_lut_11313.LUT_INIT = 16'he4aa;
    SB_LUT4 n12617_bdd_4_lut (.I0(n12617), .I1(ram_s_109_5), .I2(ram_s_108_5), 
            .I3(port_id[1]), .O(n12620));
    defparam n12617_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10855 (.I0(port_id[2]), .I1(n10481), .I2(n10499), 
            .I3(port_id[3]), .O(n12017));
    defparam port_id_2__bdd_4_lut_10855.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11308 (.I0(port_id[0]), .I1(ram_s_94_4), 
            .I2(ram_s_95_4), .I3(port_id[1]), .O(n12611));
    defparam port_id_0__bdd_4_lut_11308.LUT_INIT = 16'he4aa;
    SB_LUT4 n12611_bdd_4_lut (.I0(n12611), .I1(ram_s_93_4), .I2(ram_s_92_4), 
            .I3(port_id[1]), .O(n9737));
    defparam n12611_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11303 (.I0(port_id[0]), .I1(ram_s_10_1), 
            .I2(ram_s_11_1), .I3(port_id[1]), .O(n12605));
    defparam port_id_0__bdd_4_lut_11303.LUT_INIT = 16'he4aa;
    SB_LUT4 n12605_bdd_4_lut (.I0(n12605), .I1(ram_s_9_1), .I2(ram_s_8_1), 
            .I3(port_id[1]), .O(n12608));
    defparam n12605_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10521 (.I0(port_id[0]), .I1(ram_s_2_5), 
            .I2(ram_s_3_5), .I3(port_id[1]), .O(n11639));
    defparam port_id_0__bdd_4_lut_10521.LUT_INIT = 16'he4aa;
    SB_LUT4 n11639_bdd_4_lut (.I0(n11639), .I1(ram_s_1_5), .I2(ram_s_0_5), 
            .I3(port_id[1]), .O(n11642));
    defparam n11639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12017_bdd_4_lut (.I0(n12017), .I1(n10457), .I2(n10445), .I3(port_id[3]), 
            .O(n12020));
    defparam n12017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11298 (.I0(port_id[0]), .I1(ram_s_34_3), 
            .I2(ram_s_35_3), .I3(port_id[1]), .O(n12599));
    defparam port_id_0__bdd_4_lut_11298.LUT_INIT = 16'he4aa;
    SB_LUT4 n12599_bdd_4_lut (.I0(n12599), .I1(ram_s_33_3), .I2(ram_s_32_3), 
            .I3(port_id[1]), .O(n10844));
    defparam n12599_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11293 (.I0(port_id[0]), .I1(ram_s_186_2), 
            .I2(ram_s_187_2), .I3(port_id[1]), .O(n12593));
    defparam port_id_0__bdd_4_lut_11293.LUT_INIT = 16'he4aa;
    SB_LUT4 n12593_bdd_4_lut (.I0(n12593), .I1(ram_s_185_2), .I2(ram_s_184_2), 
            .I3(port_id[1]), .O(n12596));
    defparam n12593_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1403_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_95_3), .O(n1651));   // src/ram.vhd(68[19:45])
    defparam i1403_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_2__bdd_4_lut_11318 (.I0(port_id[2]), .I1(n9620), .I2(n9632), 
            .I3(port_id[3]), .O(n12587));
    defparam port_id_2__bdd_4_lut_11318.LUT_INIT = 16'he4aa;
    SB_LUT4 n12587_bdd_4_lut (.I0(n12587), .I1(n9614), .I2(n9599), .I3(port_id[3]), 
            .O(n12590));
    defparam n12587_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11288 (.I0(port_id[0]), .I1(ram_s_194_7), 
            .I2(ram_s_195_7), .I3(port_id[1]), .O(n12581));
    defparam port_id_0__bdd_4_lut_11288.LUT_INIT = 16'he4aa;
    SB_LUT4 n12581_bdd_4_lut (.I0(n12581), .I1(ram_s_193_7), .I2(ram_s_192_7), 
            .I3(port_id[1]), .O(n10445));
    defparam n12581_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11283 (.I0(port_id[2]), .I1(n8963), .I2(n8975), 
            .I3(port_id[3]), .O(n12575));
    defparam port_id_2__bdd_4_lut_11283.LUT_INIT = 16'he4aa;
    SB_LUT4 n12575_bdd_4_lut (.I0(n12575), .I1(n8960), .I2(n8951), .I3(port_id[3]), 
            .O(n12578));
    defparam n12575_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11278 (.I0(port_id[0]), .I1(ram_s_98_4), 
            .I2(ram_s_99_4), .I3(port_id[1]), .O(n12569));
    defparam port_id_0__bdd_4_lut_11278.LUT_INIT = 16'he4aa;
    SB_LUT4 n12569_bdd_4_lut (.I0(n12569), .I1(ram_s_97_4), .I2(ram_s_96_4), 
            .I3(port_id[1]), .O(n9740));
    defparam n12569_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_11333 (.I0(port_id[4]), .I1(n10745), .I2(n10757), 
            .I3(port_id[5]), .O(n12563));
    defparam port_id_4__bdd_4_lut_11333.LUT_INIT = 16'he4aa;
    SB_LUT4 n12563_bdd_4_lut (.I0(n12563), .I1(n10739), .I2(n10721), .I3(port_id[5]), 
            .O(n10847));
    defparam n12563_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11005 (.I0(port_id[0]), .I1(ram_s_26_1), 
            .I2(ram_s_27_1), .I3(port_id[1]), .O(n12245));
    defparam port_id_0__bdd_4_lut_11005.LUT_INIT = 16'he4aa;
    SB_LUT4 n12245_bdd_4_lut (.I0(n12245), .I1(ram_s_25_1), .I2(ram_s_24_1), 
            .I3(port_id[1]), .O(n12248));
    defparam n12245_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10496 (.I0(port_id[0]), .I1(ram_s_138_7), 
            .I2(ram_s_139_7), .I3(port_id[1]), .O(n11633));
    defparam port_id_0__bdd_4_lut_10496.LUT_INIT = 16'he4aa;
    SB_LUT4 n11633_bdd_4_lut (.I0(n11633), .I1(ram_s_137_7), .I2(ram_s_136_7), 
            .I3(port_id[1]), .O(n11636));
    defparam n11633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11000 (.I0(port_id[0]), .I1(ram_s_30_2), 
            .I2(ram_s_31_2), .I3(port_id[1]), .O(n12239));
    defparam port_id_0__bdd_4_lut_11000.LUT_INIT = 16'he4aa;
    SB_LUT4 n12239_bdd_4_lut (.I0(n12239), .I1(ram_s_29_2), .I2(ram_s_28_2), 
            .I3(port_id[1]), .O(n12242));
    defparam n12239_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11055 (.I0(port_id[2]), .I1(n8945), .I2(n8969), 
            .I3(port_id[3]), .O(n12233));
    defparam port_id_2__bdd_4_lut_11055.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_2__bdd_4_lut_10810 (.I0(port_id[2]), .I1(n9032), .I2(n9047), 
            .I3(port_id[3]), .O(n12011));
    defparam port_id_2__bdd_4_lut_10810.LUT_INIT = 16'he4aa;
    SB_LUT4 n12233_bdd_4_lut (.I0(n12233), .I1(n11954), .I2(n11354), .I3(port_id[3]), 
            .O(n12236));
    defparam n12233_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12011_bdd_4_lut (.I0(n12011), .I1(n9029), .I2(n9020), .I3(port_id[3]), 
            .O(n12014));
    defparam n12011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1402_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_95_2), .O(n1650));   // src/ram.vhd(68[19:45])
    defparam i1402_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_2__bdd_4_lut_10990 (.I0(port_id[2]), .I1(n10340), .I2(n10358), 
            .I3(port_id[3]), .O(n12227));
    defparam port_id_2__bdd_4_lut_10990.LUT_INIT = 16'he4aa;
    SB_LUT4 n12227_bdd_4_lut (.I0(n12227), .I1(n10322), .I2(n10304), .I3(port_id[3]), 
            .O(n12230));
    defparam n12227_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10645 (.I0(port_id[2]), .I1(n9188), .I2(n9200), 
            .I3(port_id[3]), .O(n11813));
    defparam port_id_2__bdd_4_lut_10645.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10491 (.I0(port_id[0]), .I1(ram_s_218_7), 
            .I2(ram_s_219_7), .I3(port_id[1]), .O(n11627));
    defparam port_id_0__bdd_4_lut_10491.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10815 (.I0(port_id[0]), .I1(ram_s_202_3), 
            .I2(ram_s_203_3), .I3(port_id[1]), .O(n12005));
    defparam port_id_0__bdd_4_lut_10815.LUT_INIT = 16'he4aa;
    SB_LUT4 n11813_bdd_4_lut (.I0(n11813), .I1(n9167), .I2(n9152), .I3(port_id[3]), 
            .O(n11816));
    defparam n11813_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12005_bdd_4_lut (.I0(n12005), .I1(ram_s_201_3), .I2(ram_s_200_3), 
            .I3(port_id[1]), .O(n12008));
    defparam n12005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_5__bdd_4_lut_11443 (.I0(port_id[5]), .I1(n11786), .I2(n8935), 
            .I3(port_id[6]), .O(n11807));
    defparam port_id_5__bdd_4_lut_11443.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10995 (.I0(port_id[0]), .I1(ram_s_102_4), 
            .I2(ram_s_103_4), .I3(port_id[1]), .O(n12221));
    defparam port_id_0__bdd_4_lut_10995.LUT_INIT = 16'he4aa;
    SB_LUT4 n11807_bdd_4_lut (.I0(n11807), .I1(n8917), .I2(n11780), .I3(port_id[6]), 
            .O(n11810));
    defparam n11807_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10805 (.I0(port_id[2]), .I1(n9368), .I2(n9395), 
            .I3(port_id[3]), .O(n11999));
    defparam port_id_2__bdd_4_lut_10805.LUT_INIT = 16'he4aa;
    SB_LUT4 n12221_bdd_4_lut (.I0(n12221), .I1(ram_s_101_4), .I2(ram_s_100_4), 
            .I3(port_id[1]), .O(n9758));
    defparam n12221_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11999_bdd_4_lut (.I0(n11999), .I1(n9323), .I2(n9302), .I3(port_id[3]), 
            .O(n12002));
    defparam n11999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut_11753 (.I0(port_id[3]), .I1(n10941), .I2(n10942), 
            .I3(port_id[4]), .O(n11801));
    defparam port_id_3__bdd_4_lut_11753.LUT_INIT = 16'he4aa;
    SB_LUT4 n11801_bdd_4_lut (.I0(n11801), .I1(n10906), .I2(n10905), .I3(port_id[4]), 
            .O(n11804));
    defparam n11801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11627_bdd_4_lut (.I0(n11627), .I1(ram_s_217_7), .I2(ram_s_216_7), 
            .I3(port_id[1]), .O(n10541));
    defparam n11627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10795 (.I0(port_id[2]), .I1(n11210), .I2(n8903), 
            .I3(port_id[3]), .O(n11993));
    defparam port_id_2__bdd_4_lut_10795.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_3__bdd_4_lut_10631 (.I0(port_id[3]), .I1(n10881), .I2(n10882), 
            .I3(port_id[4]), .O(n11795));
    defparam port_id_3__bdd_4_lut_10631.LUT_INIT = 16'he4aa;
    SB_LUT4 n11795_bdd_4_lut (.I0(n11795), .I1(n10870), .I2(n10869), .I3(port_id[4]), 
            .O(n11798));
    defparam n11795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11993_bdd_4_lut (.I0(n11993), .I1(n11282), .I2(n11312), .I3(port_id[3]), 
            .O(n11996));
    defparam n11993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10985 (.I0(port_id[2]), .I1(n9002), .I2(n9011), 
            .I3(port_id[3]), .O(n12215));
    defparam port_id_2__bdd_4_lut_10985.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11268 (.I0(port_id[0]), .I1(ram_s_90_6), 
            .I2(ram_s_91_6), .I3(port_id[1]), .O(n12557));
    defparam port_id_0__bdd_4_lut_11268.LUT_INIT = 16'he4aa;
    SB_LUT4 n12557_bdd_4_lut (.I0(n12557), .I1(ram_s_89_6), .I2(ram_s_88_6), 
            .I3(port_id[1]), .O(n12560));
    defparam n12557_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11258 (.I0(port_id[0]), .I1(ram_s_150_1), 
            .I2(ram_s_151_1), .I3(port_id[1]), .O(n12551));
    defparam port_id_0__bdd_4_lut_11258.LUT_INIT = 16'he4aa;
    SB_LUT4 n12551_bdd_4_lut (.I0(n12551), .I1(ram_s_149_1), .I2(ram_s_148_1), 
            .I3(port_id[1]), .O(n12554));
    defparam n12551_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1401_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_95_1), .O(n1649));   // src/ram.vhd(68[19:45])
    defparam i1401_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_1__bdd_4_lut_11338 (.I0(port_id[1]), .I1(n9714), .I2(n9715), 
            .I3(port_id[2]), .O(n12539));
    defparam port_id_1__bdd_4_lut_11338.LUT_INIT = 16'he4aa;
    SB_LUT4 n12539_bdd_4_lut (.I0(n12539), .I1(n9694), .I2(n9693), .I3(port_id[2]), 
            .O(n12542));
    defparam n12539_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11253 (.I0(port_id[0]), .I1(ram_s_82_7), 
            .I2(ram_s_83_7), .I3(port_id[1]), .O(n12533));
    defparam port_id_0__bdd_4_lut_11253.LUT_INIT = 16'he4aa;
    SB_LUT4 n12533_bdd_4_lut (.I0(n12533), .I1(ram_s_81_7), .I2(ram_s_80_7), 
            .I3(port_id[1]), .O(n12536));
    defparam n12533_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11273 (.I0(port_id[2]), .I1(n10088), .I2(n12494), 
            .I3(port_id[3]), .O(n12527));
    defparam port_id_2__bdd_4_lut_11273.LUT_INIT = 16'he4aa;
    SB_LUT4 n12527_bdd_4_lut (.I0(n12527), .I1(n10052), .I2(n10016), .I3(port_id[3]), 
            .O(n12530));
    defparam n12527_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11233 (.I0(port_id[2]), .I1(n10775), .I2(n10799), 
            .I3(port_id[3]), .O(n12521));
    defparam port_id_2__bdd_4_lut_11233.LUT_INIT = 16'he4aa;
    SB_LUT4 n12521_bdd_4_lut (.I0(n12521), .I1(n10730), .I2(n10709), .I3(port_id[3]), 
            .O(n12524));
    defparam n12521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12215_bdd_4_lut (.I0(n12215), .I1(n8999), .I2(n8981), .I3(port_id[3]), 
            .O(n12218));
    defparam n12215_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10486 (.I0(port_id[0]), .I1(ram_s_42_5), 
            .I2(ram_s_43_5), .I3(port_id[1]), .O(n11621));
    defparam port_id_0__bdd_4_lut_10486.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11238 (.I0(port_id[0]), .I1(ram_s_154_1), 
            .I2(ram_s_155_1), .I3(port_id[1]), .O(n12515));
    defparam port_id_0__bdd_4_lut_11238.LUT_INIT = 16'he4aa;
    SB_LUT4 n12515_bdd_4_lut (.I0(n12515), .I1(ram_s_153_1), .I2(ram_s_152_1), 
            .I3(port_id[1]), .O(n12518));
    defparam n12515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11223 (.I0(port_id[0]), .I1(ram_s_150_3), 
            .I2(ram_s_151_3), .I3(port_id[1]), .O(n12509));
    defparam port_id_0__bdd_4_lut_11223.LUT_INIT = 16'he4aa;
    SB_LUT4 n12509_bdd_4_lut (.I0(n12509), .I1(ram_s_149_3), .I2(ram_s_148_3), 
            .I3(port_id[1]), .O(n9746));
    defparam n12509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11228 (.I0(port_id[2]), .I1(n9347), .I2(n11396), 
            .I3(port_id[3]), .O(n12497));
    defparam port_id_2__bdd_4_lut_11228.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_3__bdd_4_lut_10626 (.I0(port_id[3]), .I1(n10815), .I2(n10816), 
            .I3(port_id[4]), .O(n11789));
    defparam port_id_3__bdd_4_lut_10626.LUT_INIT = 16'he4aa;
    SB_LUT4 n11789_bdd_4_lut (.I0(n11789), .I1(n10786), .I2(n10785), .I3(port_id[4]), 
            .O(n11792));
    defparam n11789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1400_3_lut_4_lut (.I0(n197), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_95_0), .O(n1648));   // src/ram.vhd(68[19:45])
    defparam i1400_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_2__bdd_4_lut_10975 (.I0(port_id[2]), .I1(n11408), .I2(n11372), 
            .I3(port_id[3]), .O(n12209));
    defparam port_id_2__bdd_4_lut_10975.LUT_INIT = 16'he4aa;
    SB_LUT4 n12209_bdd_4_lut (.I0(n12209), .I1(n11960), .I2(n11180), .I3(port_id[3]), 
            .O(n12212));
    defparam n12209_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut_10621 (.I0(port_id[3]), .I1(n10812), .I2(n10813), 
            .I3(port_id[4]), .O(n11783));
    defparam port_id_3__bdd_4_lut_10621.LUT_INIT = 16'he4aa;
    SB_LUT4 n11621_bdd_4_lut (.I0(n11621), .I1(ram_s_41_5), .I2(ram_s_40_5), 
            .I3(port_id[1]), .O(n11624));
    defparam n11621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_10456 (.I0(port_id[4]), .I1(n11054), .I2(n11072), 
            .I3(port_id[5]), .O(n11525));
    defparam port_id_4__bdd_4_lut_10456.LUT_INIT = 16'he4aa;
    SB_LUT4 n11783_bdd_4_lut (.I0(n11783), .I1(n10801), .I2(n10800), .I3(port_id[4]), 
            .O(n11786));
    defparam n11783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10800 (.I0(port_id[0]), .I1(ram_s_182_1), 
            .I2(ram_s_183_1), .I3(port_id[1]), .O(n11981));
    defparam port_id_0__bdd_4_lut_10800.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_3__bdd_4_lut_10616 (.I0(port_id[3]), .I1(n10746), .I2(n10747), 
            .I3(port_id[4]), .O(n11777));
    defparam port_id_3__bdd_4_lut_10616.LUT_INIT = 16'he4aa;
    SB_LUT4 n11777_bdd_4_lut (.I0(n11777), .I1(n10723), .I2(n10722), .I3(port_id[4]), 
            .O(n11780));
    defparam n11777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11981_bdd_4_lut (.I0(n11981), .I1(ram_s_181_1), .I2(ram_s_180_1), 
            .I3(port_id[1]), .O(n11984));
    defparam n11981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10481 (.I0(port_id[0]), .I1(ram_s_38_1), 
            .I2(ram_s_39_1), .I3(port_id[1]), .O(n11615));
    defparam port_id_0__bdd_4_lut_10481.LUT_INIT = 16'he4aa;
    SB_LUT4 n11615_bdd_4_lut (.I0(n11615), .I1(ram_s_37_1), .I2(ram_s_36_1), 
            .I3(port_id[1]), .O(n11618));
    defparam n11615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11525_bdd_4_lut (.I0(n11525), .I1(n11033), .I2(n10268), .I3(port_id[5]), 
            .O(n11528));
    defparam n11525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10685 (.I0(port_id[0]), .I1(ram_s_34_0), 
            .I2(ram_s_35_0), .I3(port_id[1]), .O(n11771));
    defparam port_id_0__bdd_4_lut_10685.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10476 (.I0(port_id[0]), .I1(ram_s_206_3), 
            .I2(ram_s_207_3), .I3(port_id[1]), .O(n11609));
    defparam port_id_0__bdd_4_lut_10476.LUT_INIT = 16'he4aa;
    SB_LUT4 n11771_bdd_4_lut (.I0(n11771), .I1(ram_s_33_0), .I2(ram_s_32_0), 
            .I3(port_id[1]), .O(n11774));
    defparam n11771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10780 (.I0(port_id[0]), .I1(ram_s_30_0), 
            .I2(ram_s_31_0), .I3(port_id[1]), .O(n11975));
    defparam port_id_0__bdd_4_lut_10780.LUT_INIT = 16'he4aa;
    SB_LUT4 n12497_bdd_4_lut (.I0(n12497), .I1(n9272), .I2(n9206), .I3(port_id[3]), 
            .O(n12500));
    defparam n12497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11218 (.I0(port_id[0]), .I1(ram_s_126_7), 
            .I2(ram_s_127_7), .I3(port_id[1]), .O(n12491));
    defparam port_id_0__bdd_4_lut_11218.LUT_INIT = 16'he4aa;
    SB_LUT4 n12491_bdd_4_lut (.I0(n12491), .I1(ram_s_125_7), .I2(ram_s_124_7), 
            .I3(port_id[1]), .O(n12494));
    defparam n12491_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2367_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_215_7), .O(n2615));   // src/ram.vhd(68[19:45])
    defparam i2367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11204 (.I0(port_id[0]), .I1(ram_s_214_5), 
            .I2(ram_s_215_5), .I3(port_id[1]), .O(n12485));
    defparam port_id_0__bdd_4_lut_11204.LUT_INIT = 16'he4aa;
    SB_LUT4 n12485_bdd_4_lut (.I0(n12485), .I1(ram_s_213_5), .I2(ram_s_212_5), 
            .I3(port_id[1]), .O(n12488));
    defparam n12485_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11199 (.I0(port_id[0]), .I1(ram_s_198_7), 
            .I2(ram_s_199_7), .I3(port_id[1]), .O(n12479));
    defparam port_id_0__bdd_4_lut_11199.LUT_INIT = 16'he4aa;
    SB_LUT4 n12479_bdd_4_lut (.I0(n12479), .I1(ram_s_197_7), .I2(ram_s_196_7), 
            .I3(port_id[1]), .O(n10457));
    defparam n12479_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_11263 (.I0(port_id[4]), .I1(n10781), .I2(n10790), 
            .I3(port_id[5]), .O(n12473));
    defparam port_id_4__bdd_4_lut_11263.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_11803 (.I0(port_id[0]), .I1(ram_s_58_4), 
            .I2(ram_s_59_4), .I3(port_id[1]), .O(n13205));
    defparam port_id_0__bdd_4_lut_11803.LUT_INIT = 16'he4aa;
    SB_LUT4 n13211_bdd_4_lut (.I0(n13211), .I1(ram_s_237_4), .I2(ram_s_236_4), 
            .I3(port_id[1]), .O(n13214));
    defparam n13211_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11818 (.I0(port_id[0]), .I1(ram_s_238_4), 
            .I2(ram_s_239_4), .I3(port_id[1]), .O(n13211));
    defparam port_id_0__bdd_4_lut_11818.LUT_INIT = 16'he4aa;
    SB_LUT4 n12473_bdd_4_lut (.I0(n12473), .I1(n10769), .I2(n10760), .I3(port_id[5]), 
            .O(n10856));
    defparam n12473_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11194 (.I0(port_id[0]), .I1(ram_s_34_5), 
            .I2(ram_s_35_5), .I3(port_id[1]), .O(n12461));
    defparam port_id_0__bdd_4_lut_11194.LUT_INIT = 16'he4aa;
    SB_LUT4 n12461_bdd_4_lut (.I0(n12461), .I1(ram_s_33_5), .I2(ram_s_32_5), 
            .I3(port_id[1]), .O(n12464));
    defparam n12461_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11209 (.I0(port_id[2]), .I1(n12164), .I2(n12044), 
            .I3(port_id[3]), .O(n12455));
    defparam port_id_2__bdd_4_lut_11209.LUT_INIT = 16'he4aa;
    SB_LUT4 n12455_bdd_4_lut (.I0(n12455), .I1(n12422), .I2(n10844), .I3(port_id[3]), 
            .O(n12458));
    defparam n12455_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_11189 (.I0(port_id[4]), .I1(n10811), .I2(n10829), 
            .I3(port_id[5]), .O(n12449));
    defparam port_id_4__bdd_4_lut_11189.LUT_INIT = 16'he4aa;
    SB_LUT4 n12449_bdd_4_lut (.I0(n12449), .I1(n10805), .I2(n10793), .I3(port_id[5]), 
            .O(n10859));
    defparam n12449_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2366_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_215_6), .O(n2614));   // src/ram.vhd(68[19:45])
    defparam i2366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_11179 (.I0(port_id[0]), .I1(ram_s_14_1), 
            .I2(ram_s_15_1), .I3(port_id[1]), .O(n12443));
    defparam port_id_0__bdd_4_lut_11179.LUT_INIT = 16'he4aa;
    SB_LUT4 n12443_bdd_4_lut (.I0(n12443), .I1(ram_s_13_1), .I2(ram_s_12_1), 
            .I3(port_id[1]), .O(n12446));
    defparam n12443_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11164 (.I0(port_id[0]), .I1(ram_s_22_2), 
            .I2(ram_s_23_2), .I3(port_id[1]), .O(n12437));
    defparam port_id_0__bdd_4_lut_11164.LUT_INIT = 16'he4aa;
    SB_LUT4 n12437_bdd_4_lut (.I0(n12437), .I1(ram_s_21_2), .I2(ram_s_20_2), 
            .I3(port_id[1]), .O(n12440));
    defparam n12437_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2548_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_238_4), .O(n2796));   // src/ram.vhd(68[19:45])
    defparam i2548_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11975_bdd_4_lut (.I0(n11975), .I1(ram_s_29_0), .I2(ram_s_28_0), 
            .I3(port_id[1]), .O(n11978));
    defparam n11975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_10790 (.I0(port_id[2]), .I1(n10691), .I2(n10700), 
            .I3(port_id[3]), .O(n11969));
    defparam port_id_2__bdd_4_lut_10790.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10980 (.I0(port_id[0]), .I1(ram_s_14_0), 
            .I2(ram_s_15_0), .I3(port_id[1]), .O(n12191));
    defparam port_id_0__bdd_4_lut_10980.LUT_INIT = 16'he4aa;
    SB_LUT4 n12191_bdd_4_lut (.I0(n12191), .I1(ram_s_13_0), .I2(ram_s_12_0), 
            .I3(port_id[1]), .O(n12194));
    defparam n12191_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_11085 (.I0(port_id[1]), .I1(n9981), .I2(n9982), 
            .I3(port_id[2]), .O(n12185));
    defparam port_id_1__bdd_4_lut_11085.LUT_INIT = 16'he4aa;
    SB_LUT4 n11969_bdd_4_lut (.I0(n11969), .I1(n10670), .I2(n10655), .I3(port_id[3]), 
            .O(n11972));
    defparam n11969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12185_bdd_4_lut (.I0(n12185), .I1(n9913), .I2(n9912), .I3(port_id[2]), 
            .O(n10906));
    defparam n12185_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10955 (.I0(port_id[0]), .I1(ram_s_134_7), 
            .I2(ram_s_135_7), .I3(port_id[1]), .O(n12179));
    defparam port_id_0__bdd_4_lut_10955.LUT_INIT = 16'he4aa;
    SB_LUT4 n12179_bdd_4_lut (.I0(n12179), .I1(ram_s_133_7), .I2(ram_s_132_7), 
            .I3(port_id[1]), .O(n12182));
    defparam n12179_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10945 (.I0(port_id[0]), .I1(ram_s_218_5), 
            .I2(ram_s_219_5), .I3(port_id[1]), .O(n12173));
    defparam port_id_0__bdd_4_lut_10945.LUT_INIT = 16'he4aa;
    SB_LUT4 n12173_bdd_4_lut (.I0(n12173), .I1(ram_s_217_5), .I2(ram_s_216_5), 
            .I3(port_id[1]), .O(n12176));
    defparam n12173_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10940 (.I0(port_id[0]), .I1(ram_s_166_1), 
            .I2(ram_s_167_1), .I3(port_id[1]), .O(n12167));
    defparam port_id_0__bdd_4_lut_10940.LUT_INIT = 16'he4aa;
    SB_LUT4 n12167_bdd_4_lut (.I0(n12167), .I1(ram_s_165_1), .I2(ram_s_164_1), 
            .I3(port_id[1]), .O(n12170));
    defparam n12167_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10935 (.I0(port_id[0]), .I1(ram_s_42_3), 
            .I2(ram_s_43_3), .I3(port_id[1]), .O(n12161));
    defparam port_id_0__bdd_4_lut_10935.LUT_INIT = 16'he4aa;
    SB_LUT4 n12161_bdd_4_lut (.I0(n12161), .I1(ram_s_41_3), .I2(ram_s_40_3), 
            .I3(port_id[1]), .O(n12164));
    defparam n12161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2365_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_215_5), .O(n2613));   // src/ram.vhd(68[19:45])
    defparam i2365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10775 (.I0(port_id[0]), .I1(ram_s_54_0), 
            .I2(ram_s_55_0), .I3(port_id[1]), .O(n11963));
    defparam port_id_0__bdd_4_lut_10775.LUT_INIT = 16'he4aa;
    SB_LUT4 n11963_bdd_4_lut (.I0(n11963), .I1(ram_s_53_0), .I2(ram_s_52_0), 
            .I3(port_id[1]), .O(n11966));
    defparam n11963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1262_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_77_6), .O(n1510));   // src/ram.vhd(68[19:45])
    defparam i1262_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_0__bdd_4_lut_10606 (.I0(port_id[0]), .I1(ram_s_186_1), 
            .I2(ram_s_187_1), .I3(port_id[1]), .O(n11765));
    defparam port_id_0__bdd_4_lut_10606.LUT_INIT = 16'he4aa;
    SB_LUT4 n11765_bdd_4_lut (.I0(n11765), .I1(ram_s_185_1), .I2(ram_s_184_1), 
            .I3(port_id[1]), .O(n11768));
    defparam n11765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2364_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_215_4), .O(n2612));   // src/ram.vhd(68[19:45])
    defparam i2364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11609_bdd_4_lut (.I0(n11609), .I1(ram_s_205_3), .I2(ram_s_204_3), 
            .I3(port_id[1]), .O(n11612));
    defparam n11609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10930 (.I0(port_id[0]), .I1(ram_s_170_1), 
            .I2(ram_s_171_1), .I3(port_id[1]), .O(n12155));
    defparam port_id_0__bdd_4_lut_10930.LUT_INIT = 16'he4aa;
    SB_LUT4 port_id_0__bdd_4_lut_10765 (.I0(port_id[0]), .I1(ram_s_54_2), 
            .I2(ram_s_55_2), .I3(port_id[1]), .O(n11957));
    defparam port_id_0__bdd_4_lut_10765.LUT_INIT = 16'he4aa;
    SB_LUT4 i2547_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_238_3), .O(n2795));   // src/ram.vhd(68[19:45])
    defparam i2547_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11957_bdd_4_lut (.I0(n11957), .I1(ram_s_53_2), .I2(ram_s_52_2), 
            .I3(port_id[1]), .O(n11960));
    defparam n11957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1250_3_lut_4_lut (.I0(n159), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_76_2), .O(n1498));   // src/ram.vhd(68[19:45])
    defparam i1250_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_1__bdd_4_lut_11243 (.I0(port_id[1]), .I1(n9987), .I2(n9988), 
            .I3(port_id[2]), .O(n12425));
    defparam port_id_1__bdd_4_lut_11243.LUT_INIT = 16'he4aa;
    SB_LUT4 n12425_bdd_4_lut (.I0(n12425), .I1(n9973), .I2(n9972), .I3(port_id[2]), 
            .O(n12428));
    defparam n12425_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11159 (.I0(port_id[0]), .I1(ram_s_38_3), 
            .I2(ram_s_39_3), .I3(port_id[1]), .O(n12419));
    defparam port_id_0__bdd_4_lut_11159.LUT_INIT = 16'he4aa;
    SB_LUT4 n12419_bdd_4_lut (.I0(n12419), .I1(ram_s_37_3), .I2(ram_s_36_3), 
            .I3(port_id[1]), .O(n12422));
    defparam n12419_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11144 (.I0(port_id[0]), .I1(ram_s_18_1), 
            .I2(ram_s_19_1), .I3(port_id[1]), .O(n12413));
    defparam port_id_0__bdd_4_lut_11144.LUT_INIT = 16'he4aa;
    SB_LUT4 n12413_bdd_4_lut (.I0(n12413), .I1(ram_s_17_1), .I2(ram_s_16_1), 
            .I3(port_id[1]), .O(n12416));
    defparam n12413_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_6__bdd_4_lut_11748 (.I0(port_id[6]), .I1(n12278), .I2(n10331), 
            .I3(port_id[7]), .O(n12407));
    defparam port_id_6__bdd_4_lut_11748.LUT_INIT = 16'he4aa;
    SB_LUT4 n12407_bdd_4_lut (.I0(n12407), .I1(n9893), .I2(n9608), .I3(port_id[7]), 
            .O(spm_ram_data[6]));
    defparam n12407_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11174 (.I0(port_id[2]), .I1(n10013), .I2(n10037), 
            .I3(port_id[3]), .O(n12401));
    defparam port_id_2__bdd_4_lut_11174.LUT_INIT = 16'he4aa;
    SB_LUT4 n12401_bdd_4_lut (.I0(n12401), .I1(n9998), .I2(n9977), .I3(port_id[3]), 
            .O(n12404));
    defparam n12401_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11139 (.I0(port_id[0]), .I1(ram_s_194_3), 
            .I2(ram_s_195_3), .I3(port_id[1]), .O(n12395));
    defparam port_id_0__bdd_4_lut_11139.LUT_INIT = 16'he4aa;
    SB_LUT4 n12395_bdd_4_lut (.I0(n12395), .I1(ram_s_193_3), .I2(ram_s_192_3), 
            .I3(port_id[1]), .O(n12398));
    defparam n12395_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2363_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_215_3), .O(n2611));   // src/ram.vhd(68[19:45])
    defparam i2363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12155_bdd_4_lut (.I0(n12155), .I1(ram_s_169_1), .I2(ram_s_168_1), 
            .I3(port_id[1]), .O(n12158));
    defparam n12155_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10760 (.I0(port_id[0]), .I1(ram_s_54_3), 
            .I2(ram_s_55_3), .I3(port_id[1]), .O(n11951));
    defparam port_id_0__bdd_4_lut_10760.LUT_INIT = 16'he4aa;
    SB_LUT4 n11951_bdd_4_lut (.I0(n11951), .I1(ram_s_53_3), .I2(ram_s_52_3), 
            .I3(port_id[1]), .O(n11954));
    defparam n11951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10925 (.I0(port_id[0]), .I1(ram_s_106_4), 
            .I2(ram_s_107_4), .I3(port_id[1]), .O(n12143));
    defparam port_id_0__bdd_4_lut_10925.LUT_INIT = 16'he4aa;
    SB_LUT4 i2362_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_215_2), .O(n2610));   // src/ram.vhd(68[19:45])
    defparam i2362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2361_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_215_1), .O(n2609));   // src/ram.vhd(68[19:45])
    defparam i2361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_0__bdd_4_lut_10471 (.I0(port_id[0]), .I1(ram_s_110_4), 
            .I2(ram_s_111_4), .I3(port_id[1]), .O(n11603));
    defparam port_id_0__bdd_4_lut_10471.LUT_INIT = 16'he4aa;
    SB_LUT4 n11603_bdd_4_lut (.I0(n11603), .I1(ram_s_109_4), .I2(ram_s_108_4), 
            .I3(port_id[1]), .O(n11606));
    defparam n11603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2360_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_215_0), .O(n2608));   // src/ram.vhd(68[19:45])
    defparam i2360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 port_id_2__bdd_4_lut_10640 (.I0(port_id[2]), .I1(n10826), .I2(n11006), 
            .I3(port_id[3]), .O(n11753));
    defparam port_id_2__bdd_4_lut_10640.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i182_2_lut_3_lut (.I0(n53), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n182_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i182_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 n12143_bdd_4_lut (.I0(n12143), .I1(ram_s_105_4), .I2(ram_s_104_4), 
            .I3(port_id[1]), .O(n9764));
    defparam n12143_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11753_bdd_4_lut (.I0(n11753), .I1(n10469), .I2(n11642), .I3(port_id[3]), 
            .O(n10529));
    defparam n11753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_10466 (.I0(port_id[0]), .I1(ram_s_114_4), 
            .I2(ram_s_115_4), .I3(port_id[1]), .O(n11597));
    defparam port_id_0__bdd_4_lut_10466.LUT_INIT = 16'he4aa;
    SB_LUT4 i2546_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_238_2), .O(n2794));   // src/ram.vhd(68[19:45])
    defparam i2546_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11597_bdd_4_lut (.I0(n11597), .I1(ram_s_113_4), .I2(ram_s_112_4), 
            .I3(port_id[1]), .O(n11600));
    defparam n11597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2545_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_238_1), .O(n2793));   // src/ram.vhd(68[19:45])
    defparam i2545_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1261_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_77_5), .O(n1509));   // src/ram.vhd(68[19:45])
    defparam i1261_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i181_2_lut_3_lut (.I0(n53), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n181));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i181_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1260_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_77_4), .O(n1508));   // src/ram.vhd(68[19:45])
    defparam i1260_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_4__bdd_4_lut_10536 (.I0(port_id[4]), .I1(n10718), .I2(n10751), 
            .I3(port_id[5]), .O(n11591));
    defparam port_id_4__bdd_4_lut_10536.LUT_INIT = 16'he4aa;
    SB_LUT4 i2544_3_lut_4_lut (.I0(n227), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_238_0), .O(n2792));   // src/ram.vhd(68[19:45])
    defparam i2544_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1399_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_94_7), .O(n1647));   // src/ram.vhd(68[19:45])
    defparam i1399_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11591_bdd_4_lut (.I0(n11591), .I1(n10682), .I2(n10661), .I3(port_id[5]), 
            .O(n11594));
    defparam n11591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1398_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_94_6), .O(n1646));   // src/ram.vhd(68[19:45])
    defparam i1398_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1397_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_94_5), .O(n1645));   // src/ram.vhd(68[19:45])
    defparam i1397_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 port_id_6__bdd_4_lut_11134 (.I0(port_id[6]), .I1(n10856), .I2(n10859), 
            .I3(port_id[7]), .O(n12383));
    defparam port_id_6__bdd_4_lut_11134.LUT_INIT = 16'he4aa;
    SB_LUT4 n12383_bdd_4_lut (.I0(n12383), .I1(n10847), .I2(n10838), .I3(port_id[7]), 
            .O(spm_ram_data[1]));
    defparam n12383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11124 (.I0(port_id[0]), .I1(ram_s_26_2), 
            .I2(ram_s_27_2), .I3(port_id[1]), .O(n12377));
    defparam port_id_0__bdd_4_lut_11124.LUT_INIT = 16'he4aa;
    SB_LUT4 n12377_bdd_4_lut (.I0(n12377), .I1(ram_s_25_2), .I2(ram_s_24_2), 
            .I3(port_id[1]), .O(n12380));
    defparam n12377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13205_bdd_4_lut (.I0(n13205), .I1(ram_s_57_4), .I2(ram_s_56_4), 
            .I3(port_id[1]), .O(n9662));
    defparam n13205_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13229_bdd_4_lut (.I0(n13229), .I1(ram_s_133_1), .I2(ram_s_132_1), 
            .I3(port_id[1]), .O(n13232));
    defparam n13229_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11823 (.I0(port_id[0]), .I1(ram_s_134_1), 
            .I2(ram_s_135_1), .I3(port_id[1]), .O(n13229));
    defparam port_id_0__bdd_4_lut_11823.LUT_INIT = 16'he4aa;
    SB_LUT4 n13235_bdd_4_lut (.I0(n13235), .I1(ram_s_185_7), .I2(ram_s_184_7), 
            .I3(port_id[1]), .O(n10412));
    defparam n13235_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11828 (.I0(port_id[0]), .I1(ram_s_186_7), 
            .I2(ram_s_187_7), .I3(port_id[1]), .O(n13235));
    defparam port_id_0__bdd_4_lut_11828.LUT_INIT = 16'he4aa;
    SB_LUT4 n13241_bdd_4_lut (.I0(n13241), .I1(ram_s_29_3), .I2(ram_s_28_3), 
            .I3(port_id[1]), .O(n10799));
    defparam n13241_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11833 (.I0(port_id[0]), .I1(ram_s_30_3), 
            .I2(ram_s_31_3), .I3(port_id[1]), .O(n13241));
    defparam port_id_0__bdd_4_lut_11833.LUT_INIT = 16'he4aa;
    SB_LUT4 n13247_bdd_4_lut (.I0(n13247), .I1(ram_s_109_2), .I2(ram_s_108_2), 
            .I3(port_id[1]), .O(n13250));
    defparam n13247_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11843 (.I0(port_id[0]), .I1(ram_s_110_2), 
            .I2(ram_s_111_2), .I3(port_id[1]), .O(n13247));
    defparam port_id_0__bdd_4_lut_11843.LUT_INIT = 16'he4aa;
    SB_LUT4 n13253_bdd_4_lut (.I0(n13253), .I1(n9454), .I2(n9453), .I3(port_id[2]), 
            .O(n13256));
    defparam n13253_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_12093 (.I0(port_id[1]), .I1(n9480), .I2(n9481), 
            .I3(port_id[2]), .O(n13253));
    defparam port_id_1__bdd_4_lut_12093.LUT_INIT = 16'he4aa;
    SB_LUT4 n13259_bdd_4_lut (.I0(n13259), .I1(ram_s_5_2), .I2(ram_s_4_2), 
            .I3(port_id[1]), .O(n10796));
    defparam n13259_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11858 (.I0(port_id[0]), .I1(ram_s_6_2), 
            .I2(ram_s_7_2), .I3(port_id[1]), .O(n13259));
    defparam port_id_0__bdd_4_lut_11858.LUT_INIT = 16'he4aa;
    SB_LUT4 i1396_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_94_4), .O(n1644));   // src/ram.vhd(68[19:45])
    defparam i1396_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13277_bdd_4_lut (.I0(n13277), .I1(ram_s_101_3), .I2(ram_s_100_3), 
            .I3(port_id[1]), .O(n9323));
    defparam n13277_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11863 (.I0(port_id[0]), .I1(ram_s_102_3), 
            .I2(ram_s_103_3), .I3(port_id[1]), .O(n13277));
    defparam port_id_0__bdd_4_lut_11863.LUT_INIT = 16'he4aa;
    SB_LUT4 n13283_bdd_4_lut (.I0(n13283), .I1(ram_s_209_5), .I2(ram_s_208_5), 
            .I3(port_id[1]), .O(n13286));
    defparam n13283_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11868 (.I0(port_id[0]), .I1(ram_s_210_5), 
            .I2(ram_s_211_5), .I3(port_id[1]), .O(n13283));
    defparam port_id_0__bdd_4_lut_11868.LUT_INIT = 16'he4aa;
    SB_LUT4 n13289_bdd_4_lut (.I0(n13289), .I1(ram_s_137_3), .I2(ram_s_136_3), 
            .I3(port_id[1]), .O(n9650));
    defparam n13289_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11873 (.I0(port_id[0]), .I1(ram_s_138_3), 
            .I2(ram_s_139_3), .I3(port_id[1]), .O(n13289));
    defparam port_id_0__bdd_4_lut_11873.LUT_INIT = 16'he4aa;
    SB_LUT4 n13295_bdd_4_lut (.I0(n13295), .I1(ram_s_173_2), .I2(ram_s_172_2), 
            .I3(port_id[1]), .O(n13298));
    defparam n13295_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11883 (.I0(port_id[0]), .I1(ram_s_174_2), 
            .I2(ram_s_175_2), .I3(port_id[1]), .O(n13295));
    defparam port_id_0__bdd_4_lut_11883.LUT_INIT = 16'he4aa;
    SB_LUT4 n13301_bdd_4_lut (.I0(n13301), .I1(n11432), .I2(n11588), .I3(port_id[3]), 
            .O(n10793));
    defparam n13301_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11928 (.I0(port_id[2]), .I1(n11222), .I2(n10577), 
            .I3(port_id[3]), .O(n13301));
    defparam port_id_2__bdd_4_lut_11928.LUT_INIT = 16'he4aa;
    SB_LUT4 n13307_bdd_4_lut (.I0(n13307), .I1(ram_s_117_7), .I2(ram_s_116_7), 
            .I3(port_id[1]), .O(n10052));
    defparam n13307_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11888 (.I0(port_id[0]), .I1(ram_s_118_7), 
            .I2(ram_s_119_7), .I3(port_id[1]), .O(n13307));
    defparam port_id_0__bdd_4_lut_11888.LUT_INIT = 16'he4aa;
    SB_LUT4 n13313_bdd_4_lut (.I0(n13313), .I1(ram_s_253_3), .I2(ram_s_252_3), 
            .I3(port_id[1]), .O(n13316));
    defparam n13313_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11893 (.I0(port_id[0]), .I1(ram_s_254_3), 
            .I2(ram_s_255_3), .I3(port_id[1]), .O(n13313));
    defparam port_id_0__bdd_4_lut_11893.LUT_INIT = 16'he4aa;
    SB_LUT4 n13319_bdd_4_lut (.I0(n13319), .I1(ram_s_69_7), .I2(ram_s_68_7), 
            .I3(port_id[1]), .O(n13322));
    defparam n13319_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11898 (.I0(port_id[0]), .I1(ram_s_70_7), 
            .I2(ram_s_71_7), .I3(port_id[1]), .O(n13319));
    defparam port_id_0__bdd_4_lut_11898.LUT_INIT = 16'he4aa;
    SB_LUT4 n13325_bdd_4_lut (.I0(n13325), .I1(ram_s_249_0), .I2(ram_s_248_0), 
            .I3(port_id[1]), .O(n13328));
    defparam n13325_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11903 (.I0(port_id[0]), .I1(ram_s_250_0), 
            .I2(ram_s_251_0), .I3(port_id[1]), .O(n13325));
    defparam port_id_0__bdd_4_lut_11903.LUT_INIT = 16'he4aa;
    SB_LUT4 n13331_bdd_4_lut (.I0(n13331), .I1(ram_s_121_0), .I2(ram_s_120_0), 
            .I3(port_id[1]), .O(n9032));
    defparam n13331_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11908 (.I0(port_id[0]), .I1(ram_s_122_0), 
            .I2(ram_s_123_0), .I3(port_id[1]), .O(n13331));
    defparam port_id_0__bdd_4_lut_11908.LUT_INIT = 16'he4aa;
    SB_LUT4 n13337_bdd_4_lut (.I0(n13337), .I1(ram_s_117_0), .I2(ram_s_116_0), 
            .I3(port_id[1]), .O(n9029));
    defparam n13337_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11913 (.I0(port_id[0]), .I1(ram_s_118_0), 
            .I2(ram_s_119_0), .I3(port_id[1]), .O(n13337));
    defparam port_id_0__bdd_4_lut_11913.LUT_INIT = 16'he4aa;
    SB_LUT4 i1395_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_94_3), .O(n1643));   // src/ram.vhd(68[19:45])
    defparam i1395_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13343_bdd_4_lut (.I0(n13343), .I1(ram_s_105_2), .I2(ram_s_104_2), 
            .I3(port_id[1]), .O(n13346));
    defparam n13343_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11918 (.I0(port_id[0]), .I1(ram_s_106_2), 
            .I2(ram_s_107_2), .I3(port_id[1]), .O(n13343));
    defparam port_id_0__bdd_4_lut_11918.LUT_INIT = 16'he4aa;
    SB_LUT4 n13349_bdd_4_lut (.I0(n13349), .I1(ram_s_53_4), .I2(ram_s_52_4), 
            .I3(port_id[1]), .O(n9644));
    defparam n13349_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11923 (.I0(port_id[0]), .I1(ram_s_54_4), 
            .I2(ram_s_55_4), .I3(port_id[1]), .O(n13349));
    defparam port_id_0__bdd_4_lut_11923.LUT_INIT = 16'he4aa;
    SB_LUT4 n13355_bdd_4_lut (.I0(n13355), .I1(ram_s_5_6), .I2(ram_s_4_6), 
            .I3(port_id[1]), .O(n9023));
    defparam n13355_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11933 (.I0(port_id[0]), .I1(ram_s_6_6), 
            .I2(ram_s_7_6), .I3(port_id[1]), .O(n13355));
    defparam port_id_0__bdd_4_lut_11933.LUT_INIT = 16'he4aa;
    SB_LUT4 n13361_bdd_4_lut (.I0(n13361), .I1(n11984), .I2(n12038), .I3(port_id[3]), 
            .O(n10790));
    defparam n13361_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11963 (.I0(port_id[2]), .I1(n11768), .I2(n11696), 
            .I3(port_id[3]), .O(n13361));
    defparam port_id_2__bdd_4_lut_11963.LUT_INIT = 16'he4aa;
    SB_LUT4 n13367_bdd_4_lut (.I0(n13367), .I1(ram_s_129_1), .I2(ram_s_128_1), 
            .I3(port_id[1]), .O(n13370));
    defparam n13367_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11938 (.I0(port_id[0]), .I1(ram_s_130_1), 
            .I2(ram_s_131_1), .I3(port_id[1]), .O(n13367));
    defparam port_id_0__bdd_4_lut_11938.LUT_INIT = 16'he4aa;
    SB_LUT4 n13373_bdd_4_lut (.I0(n13373), .I1(ram_s_233_4), .I2(ram_s_232_4), 
            .I3(port_id[1]), .O(n13376));
    defparam n13373_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11943 (.I0(port_id[0]), .I1(ram_s_234_4), 
            .I2(ram_s_235_4), .I3(port_id[1]), .O(n13373));
    defparam port_id_0__bdd_4_lut_11943.LUT_INIT = 16'he4aa;
    SB_LUT4 n13379_bdd_4_lut (.I0(n13379), .I1(ram_s_169_2), .I2(ram_s_168_2), 
            .I3(port_id[1]), .O(n13382));
    defparam n13379_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11948 (.I0(port_id[0]), .I1(ram_s_170_2), 
            .I2(ram_s_171_2), .I3(port_id[1]), .O(n13379));
    defparam port_id_0__bdd_4_lut_11948.LUT_INIT = 16'he4aa;
    SB_LUT4 n13385_bdd_4_lut (.I0(n13385), .I1(ram_s_245_2), .I2(ram_s_244_2), 
            .I3(port_id[1]), .O(n13388));
    defparam n13385_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11953 (.I0(port_id[0]), .I1(ram_s_246_2), 
            .I2(ram_s_247_2), .I3(port_id[1]), .O(n13385));
    defparam port_id_0__bdd_4_lut_11953.LUT_INIT = 16'he4aa;
    SB_LUT4 n13391_bdd_4_lut (.I0(n13391), .I1(ram_s_113_0), .I2(ram_s_112_0), 
            .I3(port_id[1]), .O(n9020));
    defparam n13391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11958 (.I0(port_id[0]), .I1(ram_s_114_0), 
            .I2(ram_s_115_0), .I3(port_id[1]), .O(n13391));
    defparam port_id_0__bdd_4_lut_11958.LUT_INIT = 16'he4aa;
    SB_LUT4 n13397_bdd_4_lut (.I0(n13397), .I1(ram_s_65_3), .I2(ram_s_64_3), 
            .I3(port_id[1]), .O(n9017));
    defparam n13397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11968 (.I0(port_id[0]), .I1(ram_s_66_3), 
            .I2(ram_s_67_3), .I3(port_id[1]), .O(n13397));
    defparam port_id_0__bdd_4_lut_11968.LUT_INIT = 16'he4aa;
    SB_LUT4 n13403_bdd_4_lut (.I0(n13403), .I1(n9509), .I2(n9479), .I3(port_id[3]), 
            .O(n13406));
    defparam n13403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_11988 (.I0(port_id[2]), .I1(n9545), .I2(n9581), 
            .I3(port_id[3]), .O(n13403));
    defparam port_id_2__bdd_4_lut_11988.LUT_INIT = 16'he4aa;
    SB_LUT4 i1394_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_94_2), .O(n1642));   // src/ram.vhd(68[19:45])
    defparam i1394_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13409_bdd_4_lut (.I0(n13409), .I1(ram_s_97_3), .I2(ram_s_96_3), 
            .I3(port_id[1]), .O(n9302));
    defparam n13409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11978 (.I0(port_id[0]), .I1(ram_s_98_3), 
            .I2(ram_s_99_3), .I3(port_id[1]), .O(n13409));
    defparam port_id_0__bdd_4_lut_11978.LUT_INIT = 16'he4aa;
    SB_LUT4 n13415_bdd_4_lut (.I0(n13415), .I1(n9932), .I2(n9911), .I3(port_id[5]), 
            .O(n10043));
    defparam n13415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12128 (.I0(port_id[4]), .I1(n9950), .I2(n9971), 
            .I3(port_id[5]), .O(n13415));
    defparam port_id_4__bdd_4_lut_12128.LUT_INIT = 16'he4aa;
    SB_LUT4 n13421_bdd_4_lut (.I0(n13421), .I1(ram_s_125_1), .I2(ram_s_124_1), 
            .I3(port_id[1]), .O(n13424));
    defparam n13421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11983 (.I0(port_id[0]), .I1(ram_s_126_1), 
            .I2(ram_s_127_1), .I3(port_id[1]), .O(n13421));
    defparam port_id_0__bdd_4_lut_11983.LUT_INIT = 16'he4aa;
    SB_LUT4 n13427_bdd_4_lut (.I0(n13427), .I1(ram_s_49_4), .I2(ram_s_48_4), 
            .I3(port_id[1]), .O(n9635));
    defparam n13427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11993 (.I0(port_id[0]), .I1(ram_s_50_4), 
            .I2(ram_s_51_4), .I3(port_id[1]), .O(n13427));
    defparam port_id_0__bdd_4_lut_11993.LUT_INIT = 16'he4aa;
    SB_LUT4 n13433_bdd_4_lut (.I0(n13433), .I1(n12170), .I2(n12266), .I3(port_id[3]), 
            .O(n10781));
    defparam n13433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12053 (.I0(port_id[2]), .I1(n12158), .I2(n12086), 
            .I3(port_id[3]), .O(n13433));
    defparam port_id_2__bdd_4_lut_12053.LUT_INIT = 16'he4aa;
    SB_LUT4 n13439_bdd_4_lut (.I0(n13439), .I1(ram_s_45_4), .I2(ram_s_44_4), 
            .I3(port_id[1]), .O(n9632));
    defparam n13439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_11998 (.I0(port_id[0]), .I1(ram_s_46_4), 
            .I2(ram_s_47_4), .I3(port_id[1]), .O(n13439));
    defparam port_id_0__bdd_4_lut_11998.LUT_INIT = 16'he4aa;
    SB_LUT4 n13445_bdd_4_lut (.I0(n13445), .I1(ram_s_29_7), .I2(ram_s_28_7), 
            .I3(port_id[1]), .O(n13448));
    defparam n13445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12003 (.I0(port_id[0]), .I1(ram_s_30_7), 
            .I2(ram_s_31_7), .I3(port_id[1]), .O(n13445));
    defparam port_id_0__bdd_4_lut_12003.LUT_INIT = 16'he4aa;
    SB_LUT4 n13451_bdd_4_lut (.I0(n13451), .I1(ram_s_229_4), .I2(ram_s_228_4), 
            .I3(port_id[1]), .O(n13454));
    defparam n13451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12013 (.I0(port_id[0]), .I1(ram_s_230_4), 
            .I2(ram_s_231_4), .I3(port_id[1]), .O(n13451));
    defparam port_id_0__bdd_4_lut_12013.LUT_INIT = 16'he4aa;
    SB_LUT4 n13457_bdd_4_lut (.I0(n13457), .I1(n11594), .I2(n11240), .I3(port_id[7]), 
            .O(spm_ram_data[5]));
    defparam n13457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_6__bdd_4_lut_12088 (.I0(port_id[6]), .I1(n8942), .I2(n8978), 
            .I3(port_id[7]), .O(n13457));
    defparam port_id_6__bdd_4_lut_12088.LUT_INIT = 16'he4aa;
    SB_LUT4 n13463_bdd_4_lut (.I0(n13463), .I1(ram_s_53_5), .I2(ram_s_52_5), 
            .I3(port_id[1]), .O(n13466));
    defparam n13463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12018 (.I0(port_id[0]), .I1(ram_s_54_5), 
            .I2(ram_s_55_5), .I3(port_id[1]), .O(n13463));
    defparam port_id_0__bdd_4_lut_12018.LUT_INIT = 16'he4aa;
    SB_LUT4 n13469_bdd_4_lut (.I0(n13469), .I1(ram_s_25_3), .I2(ram_s_24_3), 
            .I3(port_id[1]), .O(n10775));
    defparam n13469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12023 (.I0(port_id[0]), .I1(ram_s_26_3), 
            .I2(ram_s_27_3), .I3(port_id[1]), .O(n13469));
    defparam port_id_0__bdd_4_lut_12023.LUT_INIT = 16'he4aa;
    SB_LUT4 i1393_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_94_1), .O(n1641));   // src/ram.vhd(68[19:45])
    defparam i1393_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13475_bdd_4_lut (.I0(n13475), .I1(ram_s_237_0), .I2(ram_s_236_0), 
            .I3(port_id[1]), .O(n13478));
    defparam n13475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12028 (.I0(port_id[0]), .I1(ram_s_238_0), 
            .I2(ram_s_239_0), .I3(port_id[1]), .O(n13475));
    defparam port_id_0__bdd_4_lut_12028.LUT_INIT = 16'he4aa;
    SB_LUT4 n13481_bdd_4_lut (.I0(n13481), .I1(ram_s_185_5), .I2(ram_s_184_5), 
            .I3(port_id[1]), .O(n9629));
    defparam n13481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12033 (.I0(port_id[0]), .I1(ram_s_186_5), 
            .I2(ram_s_187_5), .I3(port_id[1]), .O(n13481));
    defparam port_id_0__bdd_4_lut_12033.LUT_INIT = 16'he4aa;
    SB_LUT4 n13487_bdd_4_lut (.I0(n13487), .I1(ram_s_1_2), .I2(ram_s_0_2), 
            .I3(port_id[1]), .O(n10772));
    defparam n13487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12038 (.I0(port_id[0]), .I1(ram_s_2_2), 
            .I2(ram_s_3_2), .I3(port_id[1]), .O(n13487));
    defparam port_id_0__bdd_4_lut_12038.LUT_INIT = 16'he4aa;
    SB_LUT4 n13493_bdd_4_lut (.I0(n13493), .I1(ram_s_237_6), .I2(ram_s_236_6), 
            .I3(port_id[1]), .O(n10037));
    defparam n13493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12043 (.I0(port_id[0]), .I1(ram_s_238_6), 
            .I2(ram_s_239_6), .I3(port_id[1]), .O(n13493));
    defparam port_id_0__bdd_4_lut_12043.LUT_INIT = 16'he4aa;
    SB_LUT4 n13499_bdd_4_lut (.I0(n13499), .I1(ram_s_109_0), .I2(ram_s_108_0), 
            .I3(port_id[1]), .O(n9011));
    defparam n13499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12058 (.I0(port_id[0]), .I1(ram_s_110_0), 
            .I2(ram_s_111_0), .I3(port_id[1]), .O(n13499));
    defparam port_id_0__bdd_4_lut_12058.LUT_INIT = 16'he4aa;
    SB_LUT4 n13511_bdd_4_lut (.I0(n13511), .I1(n12554), .I2(n12722), .I3(port_id[3]), 
            .O(n10769));
    defparam n13511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12068 (.I0(port_id[2]), .I1(n12518), .I2(n12320), 
            .I3(port_id[3]), .O(n13511));
    defparam port_id_2__bdd_4_lut_12068.LUT_INIT = 16'he4aa;
    SB_LUT4 n13517_bdd_4_lut (.I0(n13517), .I1(ram_s_249_3), .I2(ram_s_248_3), 
            .I3(port_id[1]), .O(n13520));
    defparam n13517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12073 (.I0(port_id[0]), .I1(ram_s_250_3), 
            .I2(ram_s_251_3), .I3(port_id[1]), .O(n13517));
    defparam port_id_0__bdd_4_lut_12073.LUT_INIT = 16'he4aa;
    SB_LUT4 n13529_bdd_4_lut (.I0(n13529), .I1(n12854), .I2(n13184), .I3(port_id[3]), 
            .O(n13532));
    defparam n13529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12103 (.I0(port_id[2]), .I1(n11726), .I2(n9437), 
            .I3(port_id[3]), .O(n13529));
    defparam port_id_2__bdd_4_lut_12103.LUT_INIT = 16'he4aa;
    SB_LUT4 n13535_bdd_4_lut (.I0(n13535), .I1(ram_s_241_2), .I2(ram_s_240_2), 
            .I3(port_id[1]), .O(n13538));
    defparam n13535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12078 (.I0(port_id[0]), .I1(ram_s_242_2), 
            .I2(ram_s_243_2), .I3(port_id[1]), .O(n13535));
    defparam port_id_0__bdd_4_lut_12078.LUT_INIT = 16'he4aa;
    SB_LUT4 i1392_3_lut_4_lut (.I0(n195_adj_858), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_94_0), .O(n1640));   // src/ram.vhd(68[19:45])
    defparam i1392_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13541_bdd_4_lut (.I0(n13541), .I1(ram_s_181_7), .I2(ram_s_180_7), 
            .I3(port_id[1]), .O(n10394));
    defparam n13541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12083 (.I0(port_id[0]), .I1(ram_s_182_7), 
            .I2(ram_s_183_7), .I3(port_id[1]), .O(n13541));
    defparam port_id_0__bdd_4_lut_12083.LUT_INIT = 16'he4aa;
    SB_LUT4 n13547_bdd_4_lut (.I0(n13547), .I1(ram_s_181_3), .I2(ram_s_180_3), 
            .I3(port_id[1]), .O(n13550));
    defparam n13547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12108 (.I0(port_id[0]), .I1(ram_s_182_3), 
            .I2(ram_s_183_3), .I3(port_id[1]), .O(n13547));
    defparam port_id_0__bdd_4_lut_12108.LUT_INIT = 16'he4aa;
    SB_LUT4 n13553_bdd_4_lut (.I0(n13553), .I1(n10706), .I2(n10697), .I3(port_id[7]), 
            .O(spm_ram_data[3]));
    defparam n13553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_6__bdd_4_lut_13237 (.I0(port_id[6]), .I1(n10727), .I2(n10742), 
            .I3(port_id[7]), .O(n13553));
    defparam port_id_6__bdd_4_lut_13237.LUT_INIT = 16'he4aa;
    SB_LUT4 n13559_bdd_4_lut (.I0(n13559), .I1(n10009), .I2(n10008), .I3(port_id[2]), 
            .O(n13562));
    defparam n13559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_12302 (.I0(port_id[1]), .I1(n10017), .I2(n10018), 
            .I3(port_id[2]), .O(n13559));
    defparam port_id_1__bdd_4_lut_12302.LUT_INIT = 16'he4aa;
    SB_LUT4 n13571_bdd_4_lut (.I0(n13571), .I1(n13232), .I2(n13370), .I3(port_id[3]), 
            .O(n10760));
    defparam n13571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12148 (.I0(port_id[2]), .I1(n12860), .I2(n12758), 
            .I3(port_id[3]), .O(n13571));
    defparam port_id_2__bdd_4_lut_12148.LUT_INIT = 16'he4aa;
    SB_LUT4 n13577_bdd_4_lut (.I0(n13577), .I1(ram_s_165_2), .I2(ram_s_164_2), 
            .I3(port_id[1]), .O(n13580));
    defparam n13577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12113 (.I0(port_id[0]), .I1(ram_s_166_2), 
            .I2(ram_s_167_2), .I3(port_id[1]), .O(n13577));
    defparam port_id_0__bdd_4_lut_12113.LUT_INIT = 16'he4aa;
    SB_LUT4 n13583_bdd_4_lut (.I0(n13583), .I1(ram_s_41_4), .I2(ram_s_40_4), 
            .I3(port_id[1]), .O(n9620));
    defparam n13583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12118 (.I0(port_id[0]), .I1(ram_s_42_4), 
            .I2(ram_s_43_4), .I3(port_id[1]), .O(n13583));
    defparam port_id_0__bdd_4_lut_12118.LUT_INIT = 16'he4aa;
    SB_LUT4 n13589_bdd_4_lut (.I0(n13589), .I1(ram_s_233_0), .I2(ram_s_232_0), 
            .I3(port_id[1]), .O(n13592));
    defparam n13589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12123 (.I0(port_id[0]), .I1(ram_s_234_0), 
            .I2(ram_s_235_0), .I3(port_id[1]), .O(n13589));
    defparam port_id_0__bdd_4_lut_12123.LUT_INIT = 16'he4aa;
    SB_LUT4 n13595_bdd_4_lut (.I0(n13595), .I1(ram_s_1_6), .I2(ram_s_0_6), 
            .I3(port_id[1]), .O(n9008));
    defparam n13595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12133 (.I0(port_id[0]), .I1(ram_s_2_6), 
            .I2(ram_s_3_6), .I3(port_id[1]), .O(n13595));
    defparam port_id_0__bdd_4_lut_12133.LUT_INIT = 16'he4aa;
    SB_LUT4 n13601_bdd_4_lut (.I0(n13601), .I1(n9866), .I2(n9836), .I3(port_id[5]), 
            .O(n10025));
    defparam n13601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12217 (.I0(port_id[4]), .I1(n9878), .I2(n9902), 
            .I3(port_id[5]), .O(n13601));
    defparam port_id_4__bdd_4_lut_12217.LUT_INIT = 16'he4aa;
    SB_LUT4 i1391_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_93_7), .O(n1639));   // src/ram.vhd(68[19:45])
    defparam i1391_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13607_bdd_4_lut (.I0(n13607), .I1(ram_s_101_2), .I2(ram_s_100_2), 
            .I3(port_id[1]), .O(n13610));
    defparam n13607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12138 (.I0(port_id[0]), .I1(ram_s_102_2), 
            .I2(ram_s_103_2), .I3(port_id[1]), .O(n13607));
    defparam port_id_0__bdd_4_lut_12138.LUT_INIT = 16'he4aa;
    SB_LUT4 n13613_bdd_4_lut (.I0(n13613), .I1(ram_s_105_0), .I2(ram_s_104_0), 
            .I3(port_id[1]), .O(n9002));
    defparam n13613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12143 (.I0(port_id[0]), .I1(ram_s_106_0), 
            .I2(ram_s_107_0), .I3(port_id[1]), .O(n13613));
    defparam port_id_0__bdd_4_lut_12143.LUT_INIT = 16'he4aa;
    SB_LUT4 n13619_bdd_4_lut (.I0(n13619), .I1(ram_s_65_7), .I2(ram_s_64_7), 
            .I3(port_id[1]), .O(n13622));
    defparam n13619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12153 (.I0(port_id[0]), .I1(ram_s_66_7), 
            .I2(ram_s_67_7), .I3(port_id[1]), .O(n13619));
    defparam port_id_0__bdd_4_lut_12153.LUT_INIT = 16'he4aa;
    SB_LUT4 n13625_bdd_4_lut (.I0(n13625), .I1(n10385), .I2(n10367), .I3(port_id[3]), 
            .O(n10757));
    defparam n13625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12188 (.I0(port_id[2]), .I1(n10391), .I2(n13424), 
            .I3(port_id[3]), .O(n13625));
    defparam port_id_2__bdd_4_lut_12188.LUT_INIT = 16'he4aa;
    SB_LUT4 n13631_bdd_4_lut (.I0(n13631), .I1(ram_s_121_1), .I2(ram_s_120_1), 
            .I3(port_id[1]), .O(n10391));
    defparam n13631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12158 (.I0(port_id[0]), .I1(ram_s_122_1), 
            .I2(ram_s_123_1), .I3(port_id[1]), .O(n13631));
    defparam port_id_0__bdd_4_lut_12158.LUT_INIT = 16'he4aa;
    SB_LUT4 n13637_bdd_4_lut (.I0(n13637), .I1(ram_s_225_4), .I2(ram_s_224_4), 
            .I3(port_id[1]), .O(n13640));
    defparam n13637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12163 (.I0(port_id[0]), .I1(ram_s_226_4), 
            .I2(ram_s_227_4), .I3(port_id[1]), .O(n13637));
    defparam port_id_0__bdd_4_lut_12163.LUT_INIT = 16'he4aa;
    SB_LUT4 n13643_bdd_4_lut (.I0(n13643), .I1(ram_s_129_5), .I2(ram_s_128_5), 
            .I3(port_id[1]), .O(n13646));
    defparam n13643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12168 (.I0(port_id[0]), .I1(ram_s_130_5), 
            .I2(ram_s_131_5), .I3(port_id[1]), .O(n13643));
    defparam port_id_0__bdd_4_lut_12168.LUT_INIT = 16'he4aa;
    SB_LUT4 n13649_bdd_4_lut (.I0(n13649), .I1(ram_s_37_4), .I2(ram_s_36_4), 
            .I3(port_id[1]), .O(n9614));
    defparam n13649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12173 (.I0(port_id[0]), .I1(ram_s_38_4), 
            .I2(ram_s_39_4), .I3(port_id[1]), .O(n13649));
    defparam port_id_0__bdd_4_lut_12173.LUT_INIT = 16'he4aa;
    SB_LUT4 n13655_bdd_4_lut (.I0(n13655), .I1(ram_s_241_5), .I2(ram_s_240_5), 
            .I3(port_id[1]), .O(n10388));
    defparam n13655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12178 (.I0(port_id[0]), .I1(ram_s_242_5), 
            .I2(ram_s_243_5), .I3(port_id[1]), .O(n13655));
    defparam port_id_0__bdd_4_lut_12178.LUT_INIT = 16'he4aa;
    SB_LUT4 n13661_bdd_4_lut (.I0(n13661), .I1(ram_s_113_7), .I2(ram_s_112_7), 
            .I3(port_id[1]), .O(n10016));
    defparam n13661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12183 (.I0(port_id[0]), .I1(ram_s_114_7), 
            .I2(ram_s_115_7), .I3(port_id[1]), .O(n13661));
    defparam port_id_0__bdd_4_lut_12183.LUT_INIT = 16'he4aa;
    SB_LUT4 n13667_bdd_4_lut (.I0(n13667), .I1(ram_s_101_0), .I2(ram_s_100_0), 
            .I3(port_id[1]), .O(n8999));
    defparam n13667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12193 (.I0(port_id[0]), .I1(ram_s_102_0), 
            .I2(ram_s_103_0), .I3(port_id[1]), .O(n13667));
    defparam port_id_0__bdd_4_lut_12193.LUT_INIT = 16'he4aa;
    SB_LUT4 i1390_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_93_6), .O(n1638));   // src/ram.vhd(68[19:45])
    defparam i1390_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13673_bdd_4_lut (.I0(n13673), .I1(n11534), .I2(n12062), .I3(port_id[3]), 
            .O(n10751));
    defparam n13673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12208 (.I0(port_id[2]), .I1(n10619), .I2(n10685), 
            .I3(port_id[3]), .O(n13673));
    defparam port_id_2__bdd_4_lut_12208.LUT_INIT = 16'he4aa;
    SB_LUT4 n13679_bdd_4_lut (.I0(n13679), .I1(ram_s_141_6), .I2(ram_s_140_6), 
            .I3(port_id[1]), .O(n13682));
    defparam n13679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12198 (.I0(port_id[0]), .I1(ram_s_142_6), 
            .I2(ram_s_143_6), .I3(port_id[1]), .O(n13679));
    defparam port_id_0__bdd_4_lut_12198.LUT_INIT = 16'he4aa;
    SB_LUT4 n13685_bdd_4_lut (.I0(n13685), .I1(ram_s_117_1), .I2(ram_s_116_1), 
            .I3(port_id[1]), .O(n10385));
    defparam n13685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12203 (.I0(port_id[0]), .I1(ram_s_118_1), 
            .I2(ram_s_119_1), .I3(port_id[1]), .O(n13685));
    defparam port_id_0__bdd_4_lut_12203.LUT_INIT = 16'he4aa;
    SB_LUT4 n13691_bdd_4_lut (.I0(n13691), .I1(ram_s_233_6), .I2(ram_s_232_6), 
            .I3(port_id[1]), .O(n10013));
    defparam n13691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12237 (.I0(port_id[0]), .I1(ram_s_234_6), 
            .I2(ram_s_235_6), .I3(port_id[1]), .O(n13691));
    defparam port_id_0__bdd_4_lut_12237.LUT_INIT = 16'he4aa;
    SB_LUT4 n13697_bdd_4_lut (.I0(n13697), .I1(n10346), .I2(n10337), .I3(port_id[3]), 
            .O(n10745));
    defparam n13697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12232 (.I0(port_id[2]), .I1(n10349), .I2(n10361), 
            .I3(port_id[3]), .O(n13697));
    defparam port_id_2__bdd_4_lut_12232.LUT_INIT = 16'he4aa;
    SB_LUT4 n13709_bdd_4_lut (.I0(n13709), .I1(n11876), .I2(n11912), .I3(port_id[5]), 
            .O(n9608));
    defparam n13709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12222 (.I0(port_id[4]), .I1(n11816), .I2(n8804), 
            .I3(port_id[5]), .O(n13709));
    defparam port_id_4__bdd_4_lut_12222.LUT_INIT = 16'he4aa;
    SB_LUT4 n13715_bdd_4_lut (.I0(n13715), .I1(n10637), .I2(n10616), .I3(port_id[5]), 
            .O(n10742));
    defparam n13715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12277 (.I0(port_id[4]), .I1(n10652), .I2(n10673), 
            .I3(port_id[5]), .O(n13715));
    defparam port_id_4__bdd_4_lut_12277.LUT_INIT = 16'he4aa;
    SB_LUT4 n13727_bdd_4_lut (.I0(n13727), .I1(n10313), .I2(n10301), .I3(port_id[3]), 
            .O(n10739));
    defparam n13727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12327 (.I0(port_id[2]), .I1(n10316), .I2(n10325), 
            .I3(port_id[3]), .O(n13727));
    defparam port_id_2__bdd_4_lut_12327.LUT_INIT = 16'he4aa;
    SB_LUT4 n13733_bdd_4_lut (.I0(n13733), .I1(ram_s_133_3), .I2(ram_s_132_3), 
            .I3(port_id[1]), .O(n9605));
    defparam n13733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12257 (.I0(port_id[0]), .I1(ram_s_134_3), 
            .I2(ram_s_135_3), .I3(port_id[1]), .O(n13733));
    defparam port_id_0__bdd_4_lut_12257.LUT_INIT = 16'he4aa;
    SB_LUT4 i1389_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_93_5), .O(n1637));   // src/ram.vhd(68[19:45])
    defparam i1389_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13757_bdd_4_lut (.I0(n13757), .I1(ram_s_177_3), .I2(ram_s_176_3), 
            .I3(port_id[1]), .O(n13760));
    defparam n13757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12262 (.I0(port_id[0]), .I1(ram_s_178_3), 
            .I2(ram_s_179_3), .I3(port_id[1]), .O(n13757));
    defparam port_id_0__bdd_4_lut_12262.LUT_INIT = 16'he4aa;
    SB_LUT4 n13763_bdd_4_lut (.I0(n13763), .I1(ram_s_237_2), .I2(ram_s_236_2), 
            .I3(port_id[1]), .O(n13766));
    defparam n13763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12267 (.I0(port_id[0]), .I1(ram_s_238_2), 
            .I2(ram_s_239_2), .I3(port_id[1]), .O(n13763));
    defparam port_id_0__bdd_4_lut_12267.LUT_INIT = 16'he4aa;
    SB_LUT4 n13769_bdd_4_lut (.I0(n13769), .I1(ram_s_21_3), .I2(ram_s_20_3), 
            .I3(port_id[1]), .O(n10730));
    defparam n13769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12272 (.I0(port_id[0]), .I1(ram_s_22_3), 
            .I2(ram_s_23_3), .I3(port_id[1]), .O(n13769));
    defparam port_id_0__bdd_4_lut_12272.LUT_INIT = 16'he4aa;
    SB_LUT4 n13775_bdd_4_lut (.I0(n13775), .I1(ram_s_105_5), .I2(ram_s_104_5), 
            .I3(port_id[1]), .O(n13778));
    defparam n13775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12287 (.I0(port_id[0]), .I1(ram_s_106_5), 
            .I2(ram_s_107_5), .I3(port_id[1]), .O(n13775));
    defparam port_id_0__bdd_4_lut_12287.LUT_INIT = 16'he4aa;
    SB_LUT4 n13781_bdd_4_lut (.I0(n13781), .I1(n11414), .I2(n11996), .I3(port_id[5]), 
            .O(n10004));
    defparam n13781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12282 (.I0(port_id[4]), .I1(n9806), .I2(n9827), 
            .I3(port_id[5]), .O(n13781));
    defparam port_id_4__bdd_4_lut_12282.LUT_INIT = 16'he4aa;
    SB_LUT4 n13787_bdd_4_lut (.I0(n13787), .I1(n11204), .I2(n11558), .I3(port_id[5]), 
            .O(n10727));
    defparam n13787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12352 (.I0(port_id[4]), .I1(n10583), .I2(n10607), 
            .I3(port_id[5]), .O(n13787));
    defparam port_id_4__bdd_4_lut_12352.LUT_INIT = 16'he4aa;
    SB_LUT4 n13793_bdd_4_lut (.I0(n13793), .I1(ram_s_33_4), .I2(ram_s_32_4), 
            .I3(port_id[1]), .O(n9599));
    defparam n13793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12292 (.I0(port_id[0]), .I1(ram_s_34_4), 
            .I2(ram_s_35_4), .I3(port_id[1]), .O(n13793));
    defparam port_id_0__bdd_4_lut_12292.LUT_INIT = 16'he4aa;
    SB_LUT4 n13799_bdd_4_lut (.I0(n13799), .I1(ram_s_245_3), .I2(ram_s_244_3), 
            .I3(port_id[1]), .O(n13802));
    defparam n13799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12297 (.I0(port_id[0]), .I1(ram_s_246_3), 
            .I2(ram_s_247_3), .I3(port_id[1]), .O(n13799));
    defparam port_id_0__bdd_4_lut_12297.LUT_INIT = 16'he4aa;
    SB_LUT4 i1388_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_93_4), .O(n1636));   // src/ram.vhd(68[19:45])
    defparam i1388_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13805_bdd_4_lut (.I0(n13805), .I1(ram_s_233_2), .I2(ram_s_232_2), 
            .I3(port_id[1]), .O(n13808));
    defparam n13805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12312 (.I0(port_id[0]), .I1(ram_s_234_2), 
            .I2(ram_s_235_2), .I3(port_id[1]), .O(n13805));
    defparam port_id_0__bdd_4_lut_12312.LUT_INIT = 16'he4aa;
    SB_LUT4 n13811_bdd_4_lut (.I0(n13811), .I1(n9133), .I2(n9132), .I3(port_id[2]), 
            .O(n13814));
    defparam n13811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_12307 (.I0(port_id[1]), .I1(n9147), .I2(n9148), 
            .I3(port_id[2]), .O(n13811));
    defparam port_id_1__bdd_4_lut_12307.LUT_INIT = 16'he4aa;
    SB_LUT4 n13817_bdd_4_lut (.I0(n13817), .I1(n9493), .I2(n9492), .I3(port_id[2]), 
            .O(n13820));
    defparam n13817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_12317 (.I0(port_id[1]), .I1(n9504), .I2(n9505), 
            .I3(port_id[2]), .O(n13817));
    defparam port_id_1__bdd_4_lut_12317.LUT_INIT = 16'he4aa;
    SB_LUT4 n13823_bdd_4_lut (.I0(n13823), .I1(ram_s_137_6), .I2(ram_s_136_6), 
            .I3(port_id[1]), .O(n13826));
    defparam n13823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12332 (.I0(port_id[0]), .I1(ram_s_138_6), 
            .I2(ram_s_139_6), .I3(port_id[1]), .O(n13823));
    defparam port_id_0__bdd_4_lut_12332.LUT_INIT = 16'he4aa;
    SB_LUT4 n13829_bdd_4_lut (.I0(n13829), .I1(n9124), .I2(n9123), .I3(port_id[2]), 
            .O(n10723));
    defparam n13829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_12347 (.I0(port_id[1]), .I1(n9156), .I2(n9157), 
            .I3(port_id[2]), .O(n13829));
    defparam port_id_1__bdd_4_lut_12347.LUT_INIT = 16'he4aa;
    SB_LUT4 n13841_bdd_4_lut (.I0(n13841), .I1(n10271), .I2(n10256), .I3(port_id[3]), 
            .O(n10721));
    defparam n13841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12362 (.I0(port_id[2]), .I1(n10277), .I2(n10295), 
            .I3(port_id[3]), .O(n13841));
    defparam port_id_2__bdd_4_lut_12362.LUT_INIT = 16'he4aa;
    SB_LUT4 n13847_bdd_4_lut (.I0(n13847), .I1(ram_s_229_6), .I2(ram_s_228_6), 
            .I3(port_id[1]), .O(n9998));
    defparam n13847_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12337 (.I0(port_id[0]), .I1(ram_s_230_6), 
            .I2(ram_s_231_6), .I3(port_id[1]), .O(n13847));
    defparam port_id_0__bdd_4_lut_12337.LUT_INIT = 16'he4aa;
    SB_LUT4 n13853_bdd_4_lut (.I0(n13853), .I1(ram_s_129_3), .I2(ram_s_128_3), 
            .I3(port_id[1]), .O(n9584));
    defparam n13853_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12342 (.I0(port_id[0]), .I1(ram_s_130_3), 
            .I2(ram_s_131_3), .I3(port_id[1]), .O(n13853));
    defparam port_id_0__bdd_4_lut_12342.LUT_INIT = 16'he4aa;
    SB_LUT4 n13859_bdd_4_lut (.I0(n13859), .I1(ram_s_165_5), .I2(ram_s_164_5), 
            .I3(port_id[1]), .O(n9272));
    defparam n13859_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12357 (.I0(port_id[0]), .I1(ram_s_166_5), 
            .I2(ram_s_167_5), .I3(port_id[1]), .O(n13859));
    defparam port_id_0__bdd_4_lut_12357.LUT_INIT = 16'he4aa;
    SB_LUT4 n13865_bdd_4_lut (.I0(n13865), .I1(n9202), .I2(n9201), .I3(port_id[2]), 
            .O(n13868));
    defparam n13865_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut_12492 (.I0(port_id[1]), .I1(n9213), .I2(n9214), 
            .I3(port_id[2]), .O(n13865));
    defparam port_id_1__bdd_4_lut_12492.LUT_INIT = 16'he4aa;
    SB_LUT4 i1387_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_93_3), .O(n1635));   // src/ram.vhd(68[19:45])
    defparam i1387_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13871_bdd_4_lut (.I0(n13871), .I1(n12692), .I2(n12908), .I3(port_id[5]), 
            .O(n9995));
    defparam n13871_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12447 (.I0(port_id[4]), .I1(n12632), .I2(n12212), 
            .I3(port_id[5]), .O(n13871));
    defparam port_id_4__bdd_4_lut_12447.LUT_INIT = 16'he4aa;
    SB_LUT4 n13877_bdd_4_lut (.I0(n13877), .I1(ram_s_61_7), .I2(ram_s_60_7), 
            .I3(port_id[1]), .O(n9581));
    defparam n13877_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12367 (.I0(port_id[0]), .I1(ram_s_62_7), 
            .I2(ram_s_63_7), .I3(port_id[1]), .O(n13877));
    defparam port_id_0__bdd_4_lut_12367.LUT_INIT = 16'he4aa;
    SB_LUT4 n13883_bdd_4_lut (.I0(n13883), .I1(n10286), .I2(n11384), .I3(port_id[3]), 
            .O(n10718));
    defparam n13883_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12372 (.I0(port_id[2]), .I1(n13778), .I2(n12620), 
            .I3(port_id[3]), .O(n13883));
    defparam port_id_2__bdd_4_lut_12372.LUT_INIT = 16'he4aa;
    SB_LUT4 n13889_bdd_4_lut (.I0(n13889), .I1(ram_s_177_7), .I2(ram_s_176_7), 
            .I3(port_id[1]), .O(n10370));
    defparam n13889_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12382 (.I0(port_id[0]), .I1(ram_s_178_7), 
            .I2(ram_s_179_7), .I3(port_id[1]), .O(n13889));
    defparam port_id_0__bdd_4_lut_12382.LUT_INIT = 16'he4aa;
    SB_LUT4 n13895_bdd_4_lut (.I0(n13895), .I1(n10229), .I2(n11270), .I3(port_id[3]), 
            .O(n10715));
    defparam n13895_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12377 (.I0(port_id[2]), .I1(n10241), .I2(n10253), 
            .I3(port_id[3]), .O(n13895));
    defparam port_id_2__bdd_4_lut_12377.LUT_INIT = 16'he4aa;
    SB_LUT4 n13901_bdd_4_lut (.I0(n13901), .I1(n11618), .I2(n12128), .I3(port_id[3]), 
            .O(n10712));
    defparam n13901_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12477 (.I0(port_id[2]), .I1(n11576), .I2(n11294), 
            .I3(port_id[3]), .O(n13901));
    defparam port_id_2__bdd_4_lut_12477.LUT_INIT = 16'he4aa;
    SB_LUT4 n13907_bdd_4_lut (.I0(n13907), .I1(ram_s_113_1), .I2(ram_s_112_1), 
            .I3(port_id[1]), .O(n10367));
    defparam n13907_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12387 (.I0(port_id[0]), .I1(ram_s_114_1), 
            .I2(ram_s_115_1), .I3(port_id[1]), .O(n13907));
    defparam port_id_0__bdd_4_lut_12387.LUT_INIT = 16'he4aa;
    SB_LUT4 n13913_bdd_4_lut (.I0(n13913), .I1(ram_s_21_4), .I2(ram_s_20_4), 
            .I3(port_id[1]), .O(n13916));
    defparam n13913_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12392 (.I0(port_id[0]), .I1(ram_s_22_4), 
            .I2(ram_s_23_4), .I3(port_id[1]), .O(n13913));
    defparam port_id_0__bdd_4_lut_12392.LUT_INIT = 16'he4aa;
    SB_LUT4 n13919_bdd_4_lut (.I0(n13919), .I1(ram_s_17_3), .I2(ram_s_16_3), 
            .I3(port_id[1]), .O(n10709));
    defparam n13919_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12397 (.I0(port_id[0]), .I1(ram_s_18_3), 
            .I2(ram_s_19_3), .I3(port_id[1]), .O(n13919));
    defparam port_id_0__bdd_4_lut_12397.LUT_INIT = 16'he4aa;
    SB_LUT4 n13925_bdd_4_lut (.I0(n13925), .I1(ram_s_89_5), .I2(ram_s_88_5), 
            .I3(port_id[1]), .O(n13928));
    defparam n13925_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12402 (.I0(port_id[0]), .I1(ram_s_90_5), 
            .I2(ram_s_91_5), .I3(port_id[1]), .O(n13925));
    defparam port_id_0__bdd_4_lut_12402.LUT_INIT = 16'he4aa;
    SB_LUT4 n13931_bdd_4_lut (.I0(n13931), .I1(ram_s_241_3), .I2(ram_s_240_3), 
            .I3(port_id[1]), .O(n13934));
    defparam n13931_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12412 (.I0(port_id[0]), .I1(ram_s_242_3), 
            .I2(ram_s_243_3), .I3(port_id[1]), .O(n13931));
    defparam port_id_0__bdd_4_lut_12412.LUT_INIT = 16'he4aa;
    SB_LUT4 i1386_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_93_2), .O(n1634));   // src/ram.vhd(68[19:45])
    defparam i1386_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13937_bdd_4_lut (.I0(n13937), .I1(n13082), .I2(n11450), .I3(port_id[4]), 
            .O(n13940));
    defparam n13937_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut_12882 (.I0(port_id[3]), .I1(n11468), .I2(n8848), 
            .I3(port_id[4]), .O(n13937));
    defparam port_id_3__bdd_4_lut_12882.LUT_INIT = 16'he4aa;
    SB_LUT4 n13943_bdd_4_lut (.I0(n13943), .I1(ram_s_161_2), .I2(ram_s_160_2), 
            .I3(port_id[1]), .O(n13946));
    defparam n13943_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12417 (.I0(port_id[0]), .I1(ram_s_162_2), 
            .I2(ram_s_163_2), .I3(port_id[1]), .O(n13943));
    defparam port_id_0__bdd_4_lut_12417.LUT_INIT = 16'he4aa;
    SB_LUT4 n13949_bdd_4_lut (.I0(n13949), .I1(ram_s_109_1), .I2(ram_s_108_1), 
            .I3(port_id[1]), .O(n10361));
    defparam n13949_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12422 (.I0(port_id[0]), .I1(ram_s_110_1), 
            .I2(ram_s_111_1), .I3(port_id[1]), .O(n13949));
    defparam port_id_0__bdd_4_lut_12422.LUT_INIT = 16'he4aa;
    SB_LUT4 n13955_bdd_4_lut (.I0(n13955), .I1(ram_s_133_6), .I2(ram_s_132_6), 
            .I3(port_id[1]), .O(n13958));
    defparam n13955_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12427 (.I0(port_id[0]), .I1(ram_s_134_6), 
            .I2(ram_s_135_6), .I3(port_id[1]), .O(n13955));
    defparam port_id_0__bdd_4_lut_12427.LUT_INIT = 16'he4aa;
    SB_LUT4 n13961_bdd_4_lut (.I0(n13961), .I1(ram_s_229_2), .I2(ram_s_228_2), 
            .I3(port_id[1]), .O(n13964));
    defparam n13961_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12432 (.I0(port_id[0]), .I1(ram_s_230_2), 
            .I2(ram_s_231_2), .I3(port_id[1]), .O(n13961));
    defparam port_id_0__bdd_4_lut_12432.LUT_INIT = 16'he4aa;
    SB_LUT4 n13967_bdd_4_lut (.I0(n13967), .I1(ram_s_109_7), .I2(ram_s_108_7), 
            .I3(port_id[1]), .O(n9980));
    defparam n13967_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12437 (.I0(port_id[0]), .I1(ram_s_110_7), 
            .I2(ram_s_111_7), .I3(port_id[1]), .O(n13967));
    defparam port_id_0__bdd_4_lut_12437.LUT_INIT = 16'he4aa;
    SB_LUT4 n13973_bdd_4_lut (.I0(n13973), .I1(ram_s_25_7), .I2(ram_s_24_7), 
            .I3(port_id[1]), .O(n13976));
    defparam n13973_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12442 (.I0(port_id[0]), .I1(ram_s_26_7), 
            .I2(ram_s_27_7), .I3(port_id[1]), .O(n13973));
    defparam port_id_0__bdd_4_lut_12442.LUT_INIT = 16'he4aa;
    SB_LUT4 n13979_bdd_4_lut (.I0(n13979), .I1(ram_s_173_7), .I2(ram_s_172_7), 
            .I3(port_id[1]), .O(n10358));
    defparam n13979_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12452 (.I0(port_id[0]), .I1(ram_s_174_7), 
            .I2(ram_s_175_7), .I3(port_id[1]), .O(n13979));
    defparam port_id_0__bdd_4_lut_12452.LUT_INIT = 16'he4aa;
    SB_LUT4 n13985_bdd_4_lut (.I0(n13985), .I1(n12074), .I2(n12116), .I3(port_id[5]), 
            .O(n10706));
    defparam n13985_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12537 (.I0(port_id[4]), .I1(n12002), .I2(n11666), 
            .I3(port_id[5]), .O(n13985));
    defparam port_id_4__bdd_4_lut_12537.LUT_INIT = 16'he4aa;
    SB_LUT4 n13991_bdd_4_lut (.I0(n13991), .I1(ram_s_225_6), .I2(ram_s_224_6), 
            .I3(port_id[1]), .O(n9977));
    defparam n13991_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12457 (.I0(port_id[0]), .I1(ram_s_226_6), 
            .I2(ram_s_227_6), .I3(port_id[1]), .O(n13991));
    defparam port_id_0__bdd_4_lut_12457.LUT_INIT = 16'he4aa;
    SB_LUT4 n13997_bdd_4_lut (.I0(n13997), .I1(ram_s_61_5), .I2(ram_s_60_5), 
            .I3(port_id[1]), .O(n14000));
    defparam n13997_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12462 (.I0(port_id[0]), .I1(ram_s_62_5), 
            .I2(ram_s_63_5), .I3(port_id[1]), .O(n13997));
    defparam port_id_0__bdd_4_lut_12462.LUT_INIT = 16'he4aa;
    SB_LUT4 i1385_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_93_1), .O(n1633));   // src/ram.vhd(68[19:45])
    defparam i1385_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14003_bdd_4_lut (.I0(n14003), .I1(ram_s_221_0), .I2(ram_s_220_0), 
            .I3(port_id[1]), .O(n14006));
    defparam n14003_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12467 (.I0(port_id[0]), .I1(ram_s_222_0), 
            .I2(ram_s_223_0), .I3(port_id[1]), .O(n14003));
    defparam port_id_0__bdd_4_lut_12467.LUT_INIT = 16'he4aa;
    SB_LUT4 n14009_bdd_4_lut (.I0(n14009), .I1(ram_s_17_4), .I2(ram_s_16_4), 
            .I3(port_id[1]), .O(n14012));
    defparam n14009_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12482 (.I0(port_id[0]), .I1(ram_s_18_4), 
            .I2(ram_s_19_4), .I3(port_id[1]), .O(n14009));
    defparam port_id_0__bdd_4_lut_12482.LUT_INIT = 16'he4aa;
    SB_LUT4 n14021_bdd_4_lut (.I0(n14021), .I1(n12302), .I2(n12416), .I3(port_id[3]), 
            .O(n10703));
    defparam n14021_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12497 (.I0(port_id[2]), .I1(n12248), .I2(n12140), 
            .I3(port_id[3]), .O(n14021));
    defparam port_id_2__bdd_4_lut_12497.LUT_INIT = 16'he4aa;
    SB_LUT4 n14027_bdd_4_lut (.I0(n14027), .I1(ram_s_149_5), .I2(ram_s_148_5), 
            .I3(port_id[1]), .O(n14030));
    defparam n14027_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12487 (.I0(port_id[0]), .I1(ram_s_150_5), 
            .I2(ram_s_151_5), .I3(port_id[1]), .O(n14027));
    defparam port_id_0__bdd_4_lut_12487.LUT_INIT = 16'he4aa;
    SB_LUT4 n14033_bdd_4_lut (.I0(n14033), .I1(ram_s_237_5), .I2(ram_s_236_5), 
            .I3(port_id[1]), .O(n10352));
    defparam n14033_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12502 (.I0(port_id[0]), .I1(ram_s_238_5), 
            .I2(ram_s_239_5), .I3(port_id[1]), .O(n14033));
    defparam port_id_0__bdd_4_lut_12502.LUT_INIT = 16'he4aa;
    SB_LUT4 n14039_bdd_4_lut (.I0(n14039), .I1(n9487), .I2(n9486), .I3(port_id[2]), 
            .O(n14042));
    defparam n14039_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_1__bdd_4_lut (.I0(port_id[1]), .I1(n9498), .I2(n9499), 
            .I3(port_id[2]), .O(n14039));
    defparam port_id_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14045_bdd_4_lut (.I0(n14045), .I1(n13388), .I2(n13538), .I3(port_id[3]), 
            .O(n9971));
    defparam n14045_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12557 (.I0(port_id[2]), .I1(n13166), .I2(n13118), 
            .I3(port_id[3]), .O(n14045));
    defparam port_id_2__bdd_4_lut_12557.LUT_INIT = 16'he4aa;
    SB_LUT4 n14051_bdd_4_lut (.I0(n14051), .I1(ram_s_93_3), .I2(ram_s_92_3), 
            .I3(port_id[1]), .O(n9251));
    defparam n14051_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12507 (.I0(port_id[0]), .I1(ram_s_94_3), 
            .I2(ram_s_95_3), .I3(port_id[1]), .O(n14051));
    defparam port_id_0__bdd_4_lut_12507.LUT_INIT = 16'he4aa;
    SB_LUT4 n14057_bdd_4_lut (.I0(n14057), .I1(ram_s_253_7), .I2(ram_s_252_7), 
            .I3(port_id[1]), .O(n10700));
    defparam n14057_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12512 (.I0(port_id[0]), .I1(ram_s_254_7), 
            .I2(ram_s_255_7), .I3(port_id[1]), .O(n14057));
    defparam port_id_0__bdd_4_lut_12512.LUT_INIT = 16'he4aa;
    SB_LUT4 n14063_bdd_4_lut (.I0(n14063), .I1(ram_s_157_2), .I2(ram_s_156_2), 
            .I3(port_id[1]), .O(n14066));
    defparam n14063_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12522 (.I0(port_id[0]), .I1(ram_s_158_2), 
            .I2(ram_s_159_2), .I3(port_id[1]), .O(n14063));
    defparam port_id_0__bdd_4_lut_12522.LUT_INIT = 16'he4aa;
    SB_LUT4 i1384_3_lut_4_lut (.I0(n193_adj_859), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_93_0), .O(n1632));   // src/ram.vhd(68[19:45])
    defparam i1384_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14075_bdd_4_lut (.I0(n14075), .I1(ram_s_105_1), .I2(ram_s_104_1), 
            .I3(port_id[1]), .O(n10349));
    defparam n14075_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12527 (.I0(port_id[0]), .I1(ram_s_106_1), 
            .I2(ram_s_107_1), .I3(port_id[1]), .O(n14075));
    defparam port_id_0__bdd_4_lut_12527.LUT_INIT = 16'he4aa;
    SB_LUT4 n14081_bdd_4_lut (.I0(n14081), .I1(ram_s_97_2), .I2(ram_s_96_2), 
            .I3(port_id[1]), .O(n14084));
    defparam n14081_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12532 (.I0(port_id[0]), .I1(ram_s_98_2), 
            .I2(ram_s_99_2), .I3(port_id[1]), .O(n14081));
    defparam port_id_0__bdd_4_lut_12532.LUT_INIT = 16'he4aa;
    SB_LUT4 n14087_bdd_4_lut (.I0(n14087), .I1(ram_s_217_0), .I2(ram_s_216_0), 
            .I3(port_id[1]), .O(n14090));
    defparam n14087_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12542 (.I0(port_id[0]), .I1(ram_s_218_0), 
            .I2(ram_s_219_0), .I3(port_id[1]), .O(n14087));
    defparam port_id_0__bdd_4_lut_12542.LUT_INIT = 16'he4aa;
    SB_LUT4 n14093_bdd_4_lut (.I0(n14093), .I1(n12524), .I2(n12806), .I3(port_id[5]), 
            .O(n10697));
    defparam n14093_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut_12702 (.I0(port_id[4]), .I1(n12458), .I2(n12236), 
            .I3(port_id[5]), .O(n14093));
    defparam port_id_4__bdd_4_lut_12702.LUT_INIT = 16'he4aa;
    SB_LUT4 n14099_bdd_4_lut (.I0(n14099), .I1(ram_s_221_6), .I2(ram_s_220_6), 
            .I3(port_id[1]), .O(n14102));
    defparam n14099_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12547 (.I0(port_id[0]), .I1(ram_s_222_6), 
            .I2(ram_s_223_6), .I3(port_id[1]), .O(n14099));
    defparam port_id_0__bdd_4_lut_12547.LUT_INIT = 16'he4aa;
    SB_LUT4 n14105_bdd_4_lut (.I0(n14105), .I1(ram_s_101_1), .I2(ram_s_100_1), 
            .I3(port_id[1]), .O(n10346));
    defparam n14105_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12552 (.I0(port_id[0]), .I1(ram_s_102_1), 
            .I2(ram_s_103_1), .I3(port_id[1]), .O(n14105));
    defparam port_id_0__bdd_4_lut_12552.LUT_INIT = 16'he4aa;
    SB_LUT4 n14111_bdd_4_lut (.I0(n14111), .I1(ram_s_153_2), .I2(ram_s_152_2), 
            .I3(port_id[1]), .O(n14114));
    defparam n14111_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12562 (.I0(port_id[0]), .I1(ram_s_154_2), 
            .I2(ram_s_155_2), .I3(port_id[1]), .O(n14111));
    defparam port_id_0__bdd_4_lut_12562.LUT_INIT = 16'he4aa;
    SB_LUT4 n14117_bdd_4_lut (.I0(n14117), .I1(n12752), .I2(n13034), .I3(port_id[3]), 
            .O(n10694));
    defparam n14117_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12647 (.I0(port_id[2]), .I1(n12608), .I2(n12446), 
            .I3(port_id[3]), .O(n14117));
    defparam port_id_2__bdd_4_lut_12647.LUT_INIT = 16'he4aa;
    SB_LUT4 n14123_bdd_4_lut (.I0(n14123), .I1(ram_s_173_3), .I2(ram_s_172_3), 
            .I3(port_id[1]), .O(n14126));
    defparam n14123_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12567 (.I0(port_id[0]), .I1(ram_s_174_3), 
            .I2(ram_s_175_3), .I3(port_id[1]), .O(n14123));
    defparam port_id_0__bdd_4_lut_12567.LUT_INIT = 16'he4aa;
    SB_LUT4 n14129_bdd_4_lut (.I0(n14129), .I1(ram_s_249_7), .I2(ram_s_248_7), 
            .I3(port_id[1]), .O(n10691));
    defparam n14129_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12577 (.I0(port_id[0]), .I1(ram_s_250_7), 
            .I2(ram_s_251_7), .I3(port_id[1]), .O(n14129));
    defparam port_id_0__bdd_4_lut_12577.LUT_INIT = 16'he4aa;
    SB_LUT4 i2359_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_214_7), .O(n2607));   // src/ram.vhd(68[19:45])
    defparam i2359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14141_bdd_4_lut (.I0(n14141), .I1(ram_s_181_5), .I2(ram_s_180_5), 
            .I3(port_id[1]), .O(n9557));
    defparam n14141_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12582 (.I0(port_id[0]), .I1(ram_s_182_5), 
            .I2(ram_s_183_5), .I3(port_id[1]), .O(n14141));
    defparam port_id_0__bdd_4_lut_12582.LUT_INIT = 16'he4aa;
    SB_LUT4 n14147_bdd_4_lut (.I0(n14147), .I1(ram_s_49_5), .I2(ram_s_48_5), 
            .I3(port_id[1]), .O(n14150));
    defparam n14147_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12587 (.I0(port_id[0]), .I1(ram_s_50_5), 
            .I2(ram_s_51_5), .I3(port_id[1]), .O(n14147));
    defparam port_id_0__bdd_4_lut_12587.LUT_INIT = 16'he4aa;
    SB_LUT4 n14153_bdd_4_lut (.I0(n14153), .I1(ram_s_225_2), .I2(ram_s_224_2), 
            .I3(port_id[1]), .O(n14156));
    defparam n14153_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12592 (.I0(port_id[0]), .I1(ram_s_226_2), 
            .I2(ram_s_227_2), .I3(port_id[1]), .O(n14153));
    defparam port_id_0__bdd_4_lut_12592.LUT_INIT = 16'he4aa;
    SB_LUT4 n14159_bdd_4_lut (.I0(n14159), .I1(ram_s_105_7), .I2(ram_s_104_7), 
            .I3(port_id[1]), .O(n9959));
    defparam n14159_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12597 (.I0(port_id[0]), .I1(ram_s_106_7), 
            .I2(ram_s_107_7), .I3(port_id[1]), .O(n14159));
    defparam port_id_0__bdd_4_lut_12597.LUT_INIT = 16'he4aa;
    SB_LUT4 n14165_bdd_4_lut (.I0(n14165), .I1(ram_s_69_5), .I2(ram_s_68_5), 
            .I3(port_id[1]), .O(n14168));
    defparam n14165_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12602 (.I0(port_id[0]), .I1(ram_s_70_5), 
            .I2(ram_s_71_5), .I3(port_id[1]), .O(n14165));
    defparam port_id_0__bdd_4_lut_12602.LUT_INIT = 16'he4aa;
    SB_LUT4 n14171_bdd_4_lut (.I0(n14171), .I1(ram_s_237_3), .I2(ram_s_236_3), 
            .I3(port_id[1]), .O(n14174));
    defparam n14171_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12607 (.I0(port_id[0]), .I1(ram_s_238_3), 
            .I2(ram_s_239_3), .I3(port_id[1]), .O(n14171));
    defparam port_id_0__bdd_4_lut_12607.LUT_INIT = 16'he4aa;
    SB_LUT4 n14177_bdd_4_lut (.I0(n14177), .I1(ram_s_125_5), .I2(ram_s_124_5), 
            .I3(port_id[1]), .O(n10685));
    defparam n14177_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12612 (.I0(port_id[0]), .I1(ram_s_126_5), 
            .I2(ram_s_127_5), .I3(port_id[1]), .O(n14177));
    defparam port_id_0__bdd_4_lut_12612.LUT_INIT = 16'he4aa;
    SB_LUT4 n14183_bdd_4_lut (.I0(n14183), .I1(ram_s_129_6), .I2(ram_s_128_6), 
            .I3(port_id[1]), .O(n14186));
    defparam n14183_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12617 (.I0(port_id[0]), .I1(ram_s_130_6), 
            .I2(ram_s_131_6), .I3(port_id[1]), .O(n14183));
    defparam port_id_0__bdd_4_lut_12617.LUT_INIT = 16'he4aa;
    SB_LUT4 n14189_bdd_4_lut (.I0(n14189), .I1(ram_s_77_2), .I2(ram_s_76_2), 
            .I3(port_id[1]), .O(n8903));
    defparam n14189_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12627 (.I0(port_id[0]), .I1(ram_s_78_2), 
            .I2(ram_s_79_2), .I3(port_id[1]), .O(n14189));
    defparam port_id_0__bdd_4_lut_12627.LUT_INIT = 16'he4aa;
    SB_LUT4 n14195_bdd_4_lut (.I0(n14195), .I1(n8953), .I2(n11798), .I3(port_id[6]), 
            .O(n14198));
    defparam n14195_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_5__bdd_4_lut_12857 (.I0(port_id[5]), .I1(n8970), .I2(n8971), 
            .I3(port_id[6]), .O(n14195));
    defparam port_id_5__bdd_4_lut_12857.LUT_INIT = 16'he4aa;
    SB_LUT4 i2358_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_214_6), .O(n2606));   // src/ram.vhd(68[19:45])
    defparam i2358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14201_bdd_4_lut (.I0(n14201), .I1(ram_s_97_0), .I2(ram_s_96_0), 
            .I3(port_id[1]), .O(n8981));
    defparam n14201_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12632 (.I0(port_id[0]), .I1(ram_s_98_0), 
            .I2(ram_s_99_0), .I3(port_id[1]), .O(n14201));
    defparam port_id_0__bdd_4_lut_12632.LUT_INIT = 16'he4aa;
    SB_LUT4 n14207_bdd_4_lut (.I0(n14207), .I1(ram_s_89_3), .I2(ram_s_88_3), 
            .I3(port_id[1]), .O(n9227));
    defparam n14207_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12637 (.I0(port_id[0]), .I1(ram_s_90_3), 
            .I2(ram_s_91_3), .I3(port_id[1]), .O(n14207));
    defparam port_id_0__bdd_4_lut_12637.LUT_INIT = 16'he4aa;
    SB_LUT4 n14213_bdd_4_lut (.I0(n14213), .I1(ram_s_21_7), .I2(ram_s_20_7), 
            .I3(port_id[1]), .O(n14216));
    defparam n14213_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12642 (.I0(port_id[0]), .I1(ram_s_22_7), 
            .I2(ram_s_23_7), .I3(port_id[1]), .O(n14213));
    defparam port_id_0__bdd_4_lut_12642.LUT_INIT = 16'he4aa;
    SB_LUT4 n14219_bdd_4_lut (.I0(n14219), .I1(ram_s_169_7), .I2(ram_s_168_7), 
            .I3(port_id[1]), .O(n10340));
    defparam n14219_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12652 (.I0(port_id[0]), .I1(ram_s_170_7), 
            .I2(ram_s_171_7), .I3(port_id[1]), .O(n14219));
    defparam port_id_0__bdd_4_lut_12652.LUT_INIT = 16'he4aa;
    SB_LUT4 n14225_bdd_4_lut (.I0(n14225), .I1(n9842), .I2(n12866), .I3(port_id[3]), 
            .O(n10682));
    defparam n14225_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12672 (.I0(port_id[2]), .I1(n13928), .I2(n12914), 
            .I3(port_id[3]), .O(n14225));
    defparam port_id_2__bdd_4_lut_12672.LUT_INIT = 16'he4aa;
    SB_LUT4 n14231_bdd_4_lut (.I0(n14231), .I1(ram_s_57_7), .I2(ram_s_56_7), 
            .I3(port_id[1]), .O(n9545));
    defparam n14231_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12657 (.I0(port_id[0]), .I1(ram_s_58_7), 
            .I2(ram_s_59_7), .I3(port_id[1]), .O(n14231));
    defparam port_id_0__bdd_4_lut_12657.LUT_INIT = 16'he4aa;
    SB_LUT4 n14237_bdd_4_lut (.I0(n14237), .I1(ram_s_189_4), .I2(ram_s_188_4), 
            .I3(port_id[1]), .O(n9953));
    defparam n14237_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12662 (.I0(port_id[0]), .I1(ram_s_190_4), 
            .I2(ram_s_191_4), .I3(port_id[1]), .O(n14237));
    defparam port_id_0__bdd_4_lut_12662.LUT_INIT = 16'he4aa;
    SB_LUT4 n14243_bdd_4_lut (.I0(n14243), .I1(ram_s_253_1), .I2(ram_s_252_1), 
            .I3(port_id[1]), .O(n10679));
    defparam n14243_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12667 (.I0(port_id[0]), .I1(ram_s_254_1), 
            .I2(ram_s_255_1), .I3(port_id[1]), .O(n14243));
    defparam port_id_0__bdd_4_lut_12667.LUT_INIT = 16'he4aa;
    SB_LUT4 n14249_bdd_4_lut (.I0(n14249), .I1(ram_s_97_1), .I2(ram_s_96_1), 
            .I3(port_id[1]), .O(n10337));
    defparam n14249_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12677 (.I0(port_id[0]), .I1(ram_s_98_1), 
            .I2(ram_s_99_1), .I3(port_id[1]), .O(n14249));
    defparam port_id_0__bdd_4_lut_12677.LUT_INIT = 16'he4aa;
    SB_LUT4 n14255_bdd_4_lut (.I0(n14255), .I1(n13964), .I2(n14156), .I3(port_id[3]), 
            .O(n9950));
    defparam n14255_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12682 (.I0(port_id[2]), .I1(n13808), .I2(n13766), 
            .I3(port_id[3]), .O(n14255));
    defparam port_id_2__bdd_4_lut_12682.LUT_INIT = 16'he4aa;
    SB_LUT4 n14261_bdd_4_lut (.I0(n14261), .I1(ram_s_5_4), .I2(ram_s_4_4), 
            .I3(port_id[1]), .O(n14264));
    defparam n14261_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12687 (.I0(port_id[0]), .I1(ram_s_6_4), 
            .I2(ram_s_7_4), .I3(port_id[1]), .O(n14261));
    defparam port_id_0__bdd_4_lut_12687.LUT_INIT = 16'he4aa;
    SB_LUT4 i2357_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_214_5), .O(n2605));   // src/ram.vhd(68[19:45])
    defparam i2357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14267_bdd_4_lut (.I0(n14267), .I1(n9860), .I2(n9833), .I3(port_id[3]), 
            .O(n14270));
    defparam n14267_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12727 (.I0(port_id[2]), .I1(n9875), .I2(n9896), 
            .I3(port_id[3]), .O(n14267));
    defparam port_id_2__bdd_4_lut_12727.LUT_INIT = 16'he4aa;
    SB_LUT4 n14273_bdd_4_lut (.I0(n14273), .I1(ram_s_125_6), .I2(ram_s_124_6), 
            .I3(port_id[1]), .O(n14276));
    defparam n14273_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12692 (.I0(port_id[0]), .I1(ram_s_126_6), 
            .I2(ram_s_127_6), .I3(port_id[1]), .O(n14273));
    defparam port_id_0__bdd_4_lut_12692.LUT_INIT = 16'he4aa;
    SB_LUT4 n14279_bdd_4_lut (.I0(n14279), .I1(ram_s_249_1), .I2(ram_s_248_1), 
            .I3(port_id[1]), .O(n10676));
    defparam n14279_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12697 (.I0(port_id[0]), .I1(ram_s_250_1), 
            .I2(ram_s_251_1), .I3(port_id[1]), .O(n14279));
    defparam port_id_0__bdd_4_lut_12697.LUT_INIT = 16'he4aa;
    SB_LUT4 n14285_bdd_4_lut (.I0(n14285), .I1(ram_s_217_6), .I2(ram_s_216_6), 
            .I3(port_id[1]), .O(n14288));
    defparam n14285_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12707 (.I0(port_id[0]), .I1(ram_s_218_6), 
            .I2(ram_s_219_6), .I3(port_id[1]), .O(n14285));
    defparam port_id_0__bdd_4_lut_12707.LUT_INIT = 16'he4aa;
    SB_LUT4 n14291_bdd_4_lut (.I0(n14291), .I1(n10598), .I2(n14270), .I3(port_id[5]), 
            .O(n10331));
    defparam n14291_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_4__bdd_4_lut (.I0(port_id[4]), .I1(n12404), .I2(n9041), 
            .I3(port_id[5]), .O(n14291));
    defparam port_id_4__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14297_bdd_4_lut (.I0(n14297), .I1(ram_s_125_3), .I2(ram_s_124_3), 
            .I3(port_id[1]), .O(n9536));
    defparam n14297_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12712 (.I0(port_id[0]), .I1(ram_s_126_3), 
            .I2(ram_s_127_3), .I3(port_id[1]), .O(n14297));
    defparam port_id_0__bdd_4_lut_12712.LUT_INIT = 16'he4aa;
    SB_LUT4 n14303_bdd_4_lut (.I0(n14303), .I1(ram_s_233_3), .I2(ram_s_232_3), 
            .I3(port_id[1]), .O(n14306));
    defparam n14303_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12717 (.I0(port_id[0]), .I1(ram_s_234_3), 
            .I2(ram_s_235_3), .I3(port_id[1]), .O(n14303));
    defparam port_id_0__bdd_4_lut_12717.LUT_INIT = 16'he4aa;
    SB_LUT4 n14309_bdd_4_lut (.I0(n14309), .I1(ram_s_221_2), .I2(ram_s_220_2), 
            .I3(port_id[1]), .O(n14312));
    defparam n14309_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12722 (.I0(port_id[0]), .I1(ram_s_222_2), 
            .I2(ram_s_223_2), .I3(port_id[1]), .O(n14309));
    defparam port_id_0__bdd_4_lut_12722.LUT_INIT = 16'he4aa;
    SB_LUT4 n14315_bdd_4_lut (.I0(n14315), .I1(ram_s_93_1), .I2(ram_s_92_1), 
            .I3(port_id[1]), .O(n10325));
    defparam n14315_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12732 (.I0(port_id[0]), .I1(ram_s_94_1), 
            .I2(ram_s_95_1), .I3(port_id[1]), .O(n14315));
    defparam port_id_0__bdd_4_lut_12732.LUT_INIT = 16'he4aa;
    SB_LUT4 n14321_bdd_4_lut (.I0(n14321), .I1(n13802), .I2(n13934), .I3(port_id[3]), 
            .O(n10673));
    defparam n14321_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12742 (.I0(port_id[2]), .I1(n13520), .I2(n13316), 
            .I3(port_id[3]), .O(n14321));
    defparam port_id_2__bdd_4_lut_12742.LUT_INIT = 16'he4aa;
    SB_LUT4 n14327_bdd_4_lut (.I0(n14327), .I1(ram_s_185_4), .I2(ram_s_184_4), 
            .I3(port_id[1]), .O(n9944));
    defparam n14327_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12737 (.I0(port_id[0]), .I1(ram_s_186_4), 
            .I2(ram_s_187_4), .I3(port_id[1]), .O(n14327));
    defparam port_id_0__bdd_4_lut_12737.LUT_INIT = 16'he4aa;
    SB_LUT4 n14333_bdd_4_lut (.I0(n14333), .I1(ram_s_93_0), .I2(ram_s_92_0), 
            .I3(port_id[1]), .O(n8975));
    defparam n14333_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12747 (.I0(port_id[0]), .I1(ram_s_94_0), 
            .I2(ram_s_95_0), .I3(port_id[1]), .O(n14333));
    defparam port_id_0__bdd_4_lut_12747.LUT_INIT = 16'he4aa;
    SB_LUT4 n14339_bdd_4_lut (.I0(n14339), .I1(n11546), .I2(n12122), .I3(port_id[3]), 
            .O(n9941));
    defparam n14339_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12822 (.I0(port_id[2]), .I1(n9803), .I2(n9821), 
            .I3(port_id[3]), .O(n14339));
    defparam port_id_2__bdd_4_lut_12822.LUT_INIT = 16'he4aa;
    SB_LUT4 n14345_bdd_4_lut (.I0(n14345), .I1(ram_s_205_0), .I2(ram_s_204_0), 
            .I3(port_id[1]), .O(n14348));
    defparam n14345_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12752 (.I0(port_id[0]), .I1(ram_s_206_0), 
            .I2(ram_s_207_0), .I3(port_id[1]), .O(n14345));
    defparam port_id_0__bdd_4_lut_12752.LUT_INIT = 16'he4aa;
    SB_LUT4 n14351_bdd_4_lut (.I0(n14351), .I1(ram_s_1_4), .I2(ram_s_0_4), 
            .I3(port_id[1]), .O(n14354));
    defparam n14351_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12757 (.I0(port_id[0]), .I1(ram_s_2_4), 
            .I2(ram_s_3_4), .I3(port_id[1]), .O(n14351));
    defparam port_id_0__bdd_4_lut_12757.LUT_INIT = 16'he4aa;
    SB_LUT4 n14357_bdd_4_lut (.I0(n14357), .I1(ram_s_245_7), .I2(ram_s_244_7), 
            .I3(port_id[1]), .O(n10670));
    defparam n14357_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12762 (.I0(port_id[0]), .I1(ram_s_246_7), 
            .I2(ram_s_247_7), .I3(port_id[1]), .O(n14357));
    defparam port_id_0__bdd_4_lut_12762.LUT_INIT = 16'he4aa;
    SB_LUT4 n14363_bdd_4_lut (.I0(n14363), .I1(ram_s_165_7), .I2(ram_s_164_7), 
            .I3(port_id[1]), .O(n10322));
    defparam n14363_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12767 (.I0(port_id[0]), .I1(ram_s_166_7), 
            .I2(ram_s_167_7), .I3(port_id[1]), .O(n14363));
    defparam port_id_0__bdd_4_lut_12767.LUT_INIT = 16'he4aa;
    SB_LUT4 n14369_bdd_4_lut (.I0(n14369), .I1(ram_s_245_1), .I2(ram_s_244_1), 
            .I3(port_id[1]), .O(n10667));
    defparam n14369_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12777 (.I0(port_id[0]), .I1(ram_s_246_1), 
            .I2(ram_s_247_1), .I3(port_id[1]), .O(n14369));
    defparam port_id_0__bdd_4_lut_12777.LUT_INIT = 16'he4aa;
    SB_LUT4 n14381_bdd_4_lut (.I0(n14381), .I1(ram_s_169_3), .I2(ram_s_168_3), 
            .I3(port_id[1]), .O(n14384));
    defparam n14381_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12782 (.I0(port_id[0]), .I1(ram_s_170_3), 
            .I2(ram_s_171_3), .I3(port_id[1]), .O(n14381));
    defparam port_id_0__bdd_4_lut_12782.LUT_INIT = 16'he4aa;
    SB_LUT4 n14387_bdd_4_lut (.I0(n14387), .I1(ram_s_233_5), .I2(ram_s_232_5), 
            .I3(port_id[1]), .O(n10319));
    defparam n14387_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12787 (.I0(port_id[0]), .I1(ram_s_234_5), 
            .I2(ram_s_235_5), .I3(port_id[1]), .O(n14387));
    defparam port_id_0__bdd_4_lut_12787.LUT_INIT = 16'he4aa;
    SB_LUT4 n14393_bdd_4_lut (.I0(n14393), .I1(ram_s_89_1), .I2(ram_s_88_1), 
            .I3(port_id[1]), .O(n10316));
    defparam n14393_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12792 (.I0(port_id[0]), .I1(ram_s_90_1), 
            .I2(ram_s_91_1), .I3(port_id[1]), .O(n14393));
    defparam port_id_0__bdd_4_lut_12792.LUT_INIT = 16'he4aa;
    SB_LUT4 i2356_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_214_4), .O(n2604));   // src/ram.vhd(68[19:45])
    defparam i2356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14399_bdd_4_lut (.I0(n14399), .I1(ram_s_13_3), .I2(ram_s_12_3), 
            .I3(port_id[1]), .O(n10664));
    defparam n14399_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12797 (.I0(port_id[0]), .I1(ram_s_14_3), 
            .I2(ram_s_15_3), .I3(port_id[1]), .O(n14399));
    defparam port_id_0__bdd_4_lut_12797.LUT_INIT = 16'he4aa;
    SB_LUT4 n14405_bdd_4_lut (.I0(n14405), .I1(ram_s_85_1), .I2(ram_s_84_1), 
            .I3(port_id[1]), .O(n10313));
    defparam n14405_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12802 (.I0(port_id[0]), .I1(ram_s_86_1), 
            .I2(ram_s_87_1), .I3(port_id[1]), .O(n14405));
    defparam port_id_0__bdd_4_lut_12802.LUT_INIT = 16'he4aa;
    SB_LUT4 n14411_bdd_4_lut (.I0(n14411), .I1(ram_s_121_6), .I2(ram_s_120_6), 
            .I3(port_id[1]), .O(n14414));
    defparam n14411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12807 (.I0(port_id[0]), .I1(ram_s_122_6), 
            .I2(ram_s_123_6), .I3(port_id[1]), .O(n14411));
    defparam port_id_0__bdd_4_lut_12807.LUT_INIT = 16'he4aa;
    SB_LUT4 n14417_bdd_4_lut (.I0(n14417), .I1(ram_s_181_4), .I2(ram_s_180_4), 
            .I3(port_id[1]), .O(n9929));
    defparam n14417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12812 (.I0(port_id[0]), .I1(ram_s_182_4), 
            .I2(ram_s_183_4), .I3(port_id[1]), .O(n14417));
    defparam port_id_0__bdd_4_lut_12812.LUT_INIT = 16'he4aa;
    SB_LUT4 n14423_bdd_4_lut (.I0(n14423), .I1(ram_s_61_3), .I2(ram_s_60_3), 
            .I3(port_id[1]), .O(n8969));
    defparam n14423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12817 (.I0(port_id[0]), .I1(ram_s_62_3), 
            .I2(ram_s_63_3), .I3(port_id[1]), .O(n14423));
    defparam port_id_0__bdd_4_lut_12817.LUT_INIT = 16'he4aa;
    SB_LUT4 n14429_bdd_4_lut (.I0(n14429), .I1(ram_s_213_6), .I2(ram_s_212_6), 
            .I3(port_id[1]), .O(n14432));
    defparam n14429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12832 (.I0(port_id[0]), .I1(ram_s_214_6), 
            .I2(ram_s_215_6), .I3(port_id[1]), .O(n14429));
    defparam port_id_0__bdd_4_lut_12832.LUT_INIT = 16'he4aa;
    SB_LUT4 n14435_bdd_4_lut (.I0(n14435), .I1(n14168), .I2(n9140), .I3(port_id[3]), 
            .O(n10661));
    defparam n14435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12957 (.I0(port_id[2]), .I1(n12740), .I2(n9515), 
            .I3(port_id[3]), .O(n14435));
    defparam port_id_2__bdd_4_lut_12957.LUT_INIT = 16'he4aa;
    SB_LUT4 n14447_bdd_4_lut (.I0(n14447), .I1(ram_s_201_0), .I2(ram_s_200_0), 
            .I3(port_id[1]), .O(n14450));
    defparam n14447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12837 (.I0(port_id[0]), .I1(ram_s_202_0), 
            .I2(ram_s_203_0), .I3(port_id[1]), .O(n14447));
    defparam port_id_0__bdd_4_lut_12837.LUT_INIT = 16'he4aa;
    SB_LUT4 n14453_bdd_4_lut (.I0(n14453), .I1(ram_s_217_2), .I2(ram_s_216_2), 
            .I3(port_id[1]), .O(n14456));
    defparam n14453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12842 (.I0(port_id[0]), .I1(ram_s_218_2), 
            .I2(ram_s_219_2), .I3(port_id[1]), .O(n14453));
    defparam port_id_0__bdd_4_lut_12842.LUT_INIT = 16'he4aa;
    SB_LUT4 n14459_bdd_4_lut (.I0(n14459), .I1(ram_s_101_7), .I2(ram_s_100_7), 
            .I3(port_id[1]), .O(n9923));
    defparam n14459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12847 (.I0(port_id[0]), .I1(ram_s_102_7), 
            .I2(ram_s_103_7), .I3(port_id[1]), .O(n14459));
    defparam port_id_0__bdd_4_lut_12847.LUT_INIT = 16'he4aa;
    SB_LUT4 n14465_bdd_4_lut (.I0(n14465), .I1(ram_s_161_5), .I2(ram_s_160_5), 
            .I3(port_id[1]), .O(n9206));
    defparam n14465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12852 (.I0(port_id[0]), .I1(ram_s_162_5), 
            .I2(ram_s_163_5), .I3(port_id[1]), .O(n14465));
    defparam port_id_0__bdd_4_lut_12852.LUT_INIT = 16'he4aa;
    SB_LUT4 i2355_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_214_3), .O(n2603));   // src/ram.vhd(68[19:45])
    defparam i2355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14471_bdd_4_lut (.I0(n14471), .I1(ram_s_177_4), .I2(ram_s_176_4), 
            .I3(port_id[1]), .O(n9920));
    defparam n14471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12862 (.I0(port_id[0]), .I1(ram_s_178_4), 
            .I2(ram_s_179_4), .I3(port_id[1]), .O(n14471));
    defparam port_id_0__bdd_4_lut_12862.LUT_INIT = 16'he4aa;
    SB_LUT4 n14477_bdd_4_lut (.I0(n14477), .I1(n9502), .I2(n9501), .I3(port_id[6]), 
            .O(n14480));
    defparam n14477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_5__bdd_4_lut (.I0(port_id[5]), .I1(n13154), .I2(n9517), 
            .I3(port_id[6]), .O(n14477));
    defparam port_id_5__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14483_bdd_4_lut (.I0(n14483), .I1(ram_s_229_3), .I2(ram_s_228_3), 
            .I3(port_id[1]), .O(n14486));
    defparam n14483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12867 (.I0(port_id[0]), .I1(ram_s_230_3), 
            .I2(ram_s_231_3), .I3(port_id[1]), .O(n14483));
    defparam port_id_0__bdd_4_lut_12867.LUT_INIT = 16'he4aa;
    SB_LUT4 n14489_bdd_4_lut (.I0(n14489), .I1(ram_s_93_2), .I2(ram_s_92_2), 
            .I3(port_id[1]), .O(n8966));
    defparam n14489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12872 (.I0(port_id[0]), .I1(ram_s_94_2), 
            .I2(ram_s_95_2), .I3(port_id[1]), .O(n14489));
    defparam port_id_0__bdd_4_lut_12872.LUT_INIT = 16'he4aa;
    SB_LUT4 n14495_bdd_4_lut (.I0(n14495), .I1(ram_s_45_6), .I2(ram_s_44_6), 
            .I3(port_id[1]), .O(n9200));
    defparam n14495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12877 (.I0(port_id[0]), .I1(ram_s_46_6), 
            .I2(ram_s_47_6), .I3(port_id[1]), .O(n14495));
    defparam port_id_0__bdd_4_lut_12877.LUT_INIT = 16'he4aa;
    SB_LUT4 n14501_bdd_4_lut (.I0(n14501), .I1(ram_s_161_7), .I2(ram_s_160_7), 
            .I3(port_id[1]), .O(n10304));
    defparam n14501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12887 (.I0(port_id[0]), .I1(ram_s_162_7), 
            .I2(ram_s_163_7), .I3(port_id[1]), .O(n14501));
    defparam port_id_0__bdd_4_lut_12887.LUT_INIT = 16'he4aa;
    SB_LUT4 n14507_bdd_4_lut (.I0(n14507), .I1(n9472), .I2(n13046), .I3(port_id[4]), 
            .O(n9517));
    defparam n14507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut_13032 (.I0(port_id[3]), .I1(n13058), .I2(n9475), 
            .I3(port_id[4]), .O(n14507));
    defparam port_id_3__bdd_4_lut_13032.LUT_INIT = 16'he4aa;
    SB_LUT4 n14513_bdd_4_lut (.I0(n14513), .I1(ram_s_81_1), .I2(ram_s_80_1), 
            .I3(port_id[1]), .O(n10301));
    defparam n14513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12892 (.I0(port_id[0]), .I1(ram_s_82_1), 
            .I2(ram_s_83_1), .I3(port_id[1]), .O(n14513));
    defparam port_id_0__bdd_4_lut_12892.LUT_INIT = 16'he4aa;
    SB_LUT4 n14519_bdd_4_lut (.I0(n14519), .I1(ram_s_241_1), .I2(ram_s_240_1), 
            .I3(port_id[1]), .O(n10658));
    defparam n14519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12897 (.I0(port_id[0]), .I1(ram_s_242_1), 
            .I2(ram_s_243_1), .I3(port_id[1]), .O(n14519));
    defparam port_id_0__bdd_4_lut_12897.LUT_INIT = 16'he4aa;
    SB_LUT4 n14525_bdd_4_lut (.I0(n14525), .I1(ram_s_17_7), .I2(ram_s_16_7), 
            .I3(port_id[1]), .O(n14528));
    defparam n14525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12902 (.I0(port_id[0]), .I1(ram_s_18_7), 
            .I2(ram_s_19_7), .I3(port_id[1]), .O(n14525));
    defparam port_id_0__bdd_4_lut_12902.LUT_INIT = 16'he4aa;
    SB_LUT4 n14531_bdd_4_lut (.I0(n14531), .I1(ram_s_77_5), .I2(ram_s_76_5), 
            .I3(port_id[1]), .O(n9515));
    defparam n14531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12907 (.I0(port_id[0]), .I1(ram_s_78_5), 
            .I2(ram_s_79_5), .I3(port_id[1]), .O(n14531));
    defparam port_id_0__bdd_4_lut_12907.LUT_INIT = 16'he4aa;
    SB_LUT4 n14537_bdd_4_lut (.I0(n14537), .I1(ram_s_173_4), .I2(ram_s_172_4), 
            .I3(port_id[1]), .O(n9917));
    defparam n14537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12912 (.I0(port_id[0]), .I1(ram_s_174_4), 
            .I2(ram_s_175_4), .I3(port_id[1]), .O(n14537));
    defparam port_id_0__bdd_4_lut_12912.LUT_INIT = 16'he4aa;
    SB_LUT4 i2354_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_214_2), .O(n2602));   // src/ram.vhd(68[19:45])
    defparam i2354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14543_bdd_4_lut (.I0(n14543), .I1(ram_s_89_0), .I2(ram_s_88_0), 
            .I3(port_id[1]), .O(n8963));
    defparam n14543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12917 (.I0(port_id[0]), .I1(ram_s_90_0), 
            .I2(ram_s_91_0), .I3(port_id[1]), .O(n14543));
    defparam port_id_0__bdd_4_lut_12917.LUT_INIT = 16'he4aa;
    SB_LUT4 n14549_bdd_4_lut (.I0(n14549), .I1(ram_s_189_0), .I2(ram_s_188_0), 
            .I3(port_id[1]), .O(n14552));
    defparam n14549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12922 (.I0(port_id[0]), .I1(ram_s_190_0), 
            .I2(ram_s_191_0), .I3(port_id[1]), .O(n14549));
    defparam port_id_0__bdd_4_lut_12922.LUT_INIT = 16'he4aa;
    SB_LUT4 n14555_bdd_4_lut (.I0(n14555), .I1(ram_s_85_0), .I2(ram_s_84_0), 
            .I3(port_id[1]), .O(n8960));
    defparam n14555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12927 (.I0(port_id[0]), .I1(ram_s_86_0), 
            .I2(ram_s_87_0), .I3(port_id[1]), .O(n14555));
    defparam port_id_0__bdd_4_lut_12927.LUT_INIT = 16'he4aa;
    SB_LUT4 n14561_bdd_4_lut (.I0(n14561), .I1(ram_s_41_6), .I2(ram_s_40_6), 
            .I3(port_id[1]), .O(n9188));
    defparam n14561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12932 (.I0(port_id[0]), .I1(ram_s_42_6), 
            .I2(ram_s_43_6), .I3(port_id[1]), .O(n14561));
    defparam port_id_0__bdd_4_lut_12932.LUT_INIT = 16'he4aa;
    SB_LUT4 n14567_bdd_4_lut (.I0(n14567), .I1(ram_s_241_7), .I2(ram_s_240_7), 
            .I3(port_id[1]), .O(n10655));
    defparam n14567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12937 (.I0(port_id[0]), .I1(ram_s_242_7), 
            .I2(ram_s_243_7), .I3(port_id[1]), .O(n14567));
    defparam port_id_0__bdd_4_lut_12937.LUT_INIT = 16'he4aa;
    SB_LUT4 n14573_bdd_4_lut (.I0(n14573), .I1(ram_s_121_3), .I2(ram_s_120_3), 
            .I3(port_id[1]), .O(n9512));
    defparam n14573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12947 (.I0(port_id[0]), .I1(ram_s_122_3), 
            .I2(ram_s_123_3), .I3(port_id[1]), .O(n14573));
    defparam port_id_0__bdd_4_lut_12947.LUT_INIT = 16'he4aa;
    SB_LUT4 n14585_bdd_4_lut (.I0(n14585), .I1(ram_s_85_3), .I2(ram_s_84_3), 
            .I3(port_id[1]), .O(n9182));
    defparam n14585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12952 (.I0(port_id[0]), .I1(ram_s_86_3), 
            .I2(ram_s_87_3), .I3(port_id[1]), .O(n14585));
    defparam port_id_0__bdd_4_lut_12952.LUT_INIT = 16'he4aa;
    SB_LUT4 n14591_bdd_4_lut (.I0(n14591), .I1(ram_s_225_3), .I2(ram_s_224_3), 
            .I3(port_id[1]), .O(n14594));
    defparam n14591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12967 (.I0(port_id[0]), .I1(ram_s_226_3), 
            .I2(ram_s_227_3), .I3(port_id[1]), .O(n14591));
    defparam port_id_0__bdd_4_lut_12967.LUT_INIT = 16'he4aa;
    SB_LUT4 n14597_bdd_4_lut (.I0(n14597), .I1(n9428), .I2(n11426), .I3(port_id[3]), 
            .O(n9911));
    defparam n14597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12962 (.I0(port_id[2]), .I1(n9449), .I2(n9458), 
            .I3(port_id[3]), .O(n14597));
    defparam port_id_2__bdd_4_lut_12962.LUT_INIT = 16'he4aa;
    SB_LUT4 n14603_bdd_4_lut (.I0(n14603), .I1(n14486), .I2(n14594), .I3(port_id[3]), 
            .O(n10652));
    defparam n14603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12992 (.I0(port_id[2]), .I1(n14306), .I2(n14174), 
            .I3(port_id[3]), .O(n14603));
    defparam port_id_2__bdd_4_lut_12992.LUT_INIT = 16'he4aa;
    SB_LUT4 n14609_bdd_4_lut (.I0(n14609), .I1(ram_s_141_2), .I2(ram_s_140_2), 
            .I3(port_id[1]), .O(n14612));
    defparam n14609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12972 (.I0(port_id[0]), .I1(ram_s_142_2), 
            .I2(ram_s_143_2), .I3(port_id[1]), .O(n14609));
    defparam port_id_0__bdd_4_lut_12972.LUT_INIT = 16'he4aa;
    SB_LUT4 i2353_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_214_1), .O(n2601));   // src/ram.vhd(68[19:45])
    defparam i2353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14615_bdd_4_lut (.I0(n14615), .I1(ram_s_53_7), .I2(ram_s_52_7), 
            .I3(port_id[1]), .O(n9509));
    defparam n14615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12977 (.I0(port_id[0]), .I1(ram_s_54_7), 
            .I2(ram_s_55_7), .I3(port_id[1]), .O(n14615));
    defparam port_id_0__bdd_4_lut_12977.LUT_INIT = 16'he4aa;
    SB_LUT4 n14621_bdd_4_lut (.I0(n14621), .I1(ram_s_209_6), .I2(ram_s_208_6), 
            .I3(port_id[1]), .O(n14624));
    defparam n14621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12982 (.I0(port_id[0]), .I1(ram_s_210_6), 
            .I2(ram_s_211_6), .I3(port_id[1]), .O(n14621));
    defparam port_id_0__bdd_4_lut_12982.LUT_INIT = 16'he4aa;
    SB_LUT4 n14627_bdd_4_lut (.I0(n14627), .I1(ram_s_169_4), .I2(ram_s_168_4), 
            .I3(port_id[1]), .O(n9905));
    defparam n14627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_12987 (.I0(port_id[0]), .I1(ram_s_170_4), 
            .I2(ram_s_171_4), .I3(port_id[1]), .O(n14627));
    defparam port_id_0__bdd_4_lut_12987.LUT_INIT = 16'he4aa;
    SB_LUT4 n14633_bdd_4_lut (.I0(n14633), .I1(ram_s_237_1), .I2(ram_s_236_1), 
            .I3(port_id[1]), .O(n10649));
    defparam n14633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13007 (.I0(port_id[0]), .I1(ram_s_238_1), 
            .I2(ram_s_239_1), .I3(port_id[1]), .O(n14633));
    defparam port_id_0__bdd_4_lut_13007.LUT_INIT = 16'he4aa;
    SB_LUT4 n14639_bdd_4_lut (.I0(n14639), .I1(n13958), .I2(n14186), .I3(port_id[3]), 
            .O(n10646));
    defparam n14639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_12997 (.I0(port_id[2]), .I1(n13826), .I2(n13682), 
            .I3(port_id[3]), .O(n14639));
    defparam port_id_2__bdd_4_lut_12997.LUT_INIT = 16'he4aa;
    SB_LUT4 n14645_bdd_4_lut (.I0(n14645), .I1(n12932), .I2(n13088), .I3(port_id[3]), 
            .O(n9902));
    defparam n14645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13057 (.I0(port_id[2]), .I1(n12596), .I2(n12332), 
            .I3(port_id[3]), .O(n14645));
    defparam port_id_2__bdd_4_lut_13057.LUT_INIT = 16'he4aa;
    SB_LUT4 n14657_bdd_4_lut (.I0(n14657), .I1(ram_s_77_1), .I2(ram_s_76_1), 
            .I3(port_id[1]), .O(n10295));
    defparam n14657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13012 (.I0(port_id[0]), .I1(ram_s_78_1), 
            .I2(ram_s_79_1), .I3(port_id[1]), .O(n14657));
    defparam port_id_0__bdd_4_lut_13012.LUT_INIT = 16'he4aa;
    SB_LUT4 n14663_bdd_4_lut (.I0(n14663), .I1(ram_s_165_4), .I2(ram_s_164_4), 
            .I3(port_id[1]), .O(n9899));
    defparam n14663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13017 (.I0(port_id[0]), .I1(ram_s_166_4), 
            .I2(ram_s_167_4), .I3(port_id[1]), .O(n14663));
    defparam port_id_0__bdd_4_lut_13017.LUT_INIT = 16'he4aa;
    SB_LUT4 n14669_bdd_4_lut (.I0(n14669), .I1(ram_s_9_3), .I2(ram_s_8_3), 
            .I3(port_id[1]), .O(n10640));
    defparam n14669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13022 (.I0(port_id[0]), .I1(ram_s_10_3), 
            .I2(ram_s_11_3), .I3(port_id[1]), .O(n14669));
    defparam port_id_0__bdd_4_lut_13022.LUT_INIT = 16'he4aa;
    SB_LUT4 n14675_bdd_4_lut (.I0(n14675), .I1(ram_s_205_6), .I2(ram_s_204_6), 
            .I3(port_id[1]), .O(n9896));
    defparam n14675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13027 (.I0(port_id[0]), .I1(ram_s_206_6), 
            .I2(ram_s_207_6), .I3(port_id[1]), .O(n14675));
    defparam port_id_0__bdd_4_lut_13027.LUT_INIT = 16'he4aa;
    SB_LUT4 n14681_bdd_4_lut (.I0(n14681), .I1(ram_s_185_0), .I2(ram_s_184_0), 
            .I3(port_id[1]), .O(n14684));
    defparam n14681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13042 (.I0(port_id[0]), .I1(ram_s_186_0), 
            .I2(ram_s_187_0), .I3(port_id[1]), .O(n14681));
    defparam port_id_0__bdd_4_lut_13042.LUT_INIT = 16'he4aa;
    SB_LUT4 i2352_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_214_0), .O(n2600));   // src/ram.vhd(68[19:45])
    defparam i2352_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14687_bdd_4_lut (.I0(n14687), .I1(n13256), .I2(n11336), .I3(port_id[4]), 
            .O(n14690));
    defparam n14687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut_13037 (.I0(port_id[3]), .I1(n13820), .I2(n9847), 
            .I3(port_id[4]), .O(n14687));
    defparam port_id_3__bdd_4_lut_13037.LUT_INIT = 16'he4aa;
    SB_LUT4 n14693_bdd_4_lut (.I0(n14693), .I1(n9430), .I2(n12938), .I3(port_id[4]), 
            .O(n9502));
    defparam n14693_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_3__bdd_4_lut (.I0(port_id[3]), .I1(n12962), .I2(n9433), 
            .I3(port_id[4]), .O(n14693));
    defparam port_id_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14699_bdd_4_lut (.I0(n14699), .I1(ram_s_165_3), .I2(ram_s_164_3), 
            .I3(port_id[1]), .O(n14702));
    defparam n14699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13047 (.I0(port_id[0]), .I1(ram_s_166_3), 
            .I2(ram_s_167_3), .I3(port_id[1]), .O(n14699));
    defparam port_id_0__bdd_4_lut_13047.LUT_INIT = 16'he4aa;
    SB_LUT4 n14705_bdd_4_lut (.I0(n14705), .I1(ram_s_137_2), .I2(ram_s_136_2), 
            .I3(port_id[1]), .O(n14708));
    defparam n14705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13052 (.I0(port_id[0]), .I1(ram_s_138_2), 
            .I2(ram_s_139_2), .I3(port_id[1]), .O(n14705));
    defparam port_id_0__bdd_4_lut_13052.LUT_INIT = 16'he4aa;
    SB_LUT4 n14711_bdd_4_lut (.I0(n14711), .I1(ram_s_97_7), .I2(ram_s_96_7), 
            .I3(port_id[1]), .O(n9887));
    defparam n14711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13062 (.I0(port_id[0]), .I1(ram_s_98_7), 
            .I2(ram_s_99_7), .I3(port_id[1]), .O(n14711));
    defparam port_id_0__bdd_4_lut_13062.LUT_INIT = 16'he4aa;
    SB_LUT4 n14717_bdd_4_lut (.I0(n14717), .I1(n10232), .I2(n11228), .I3(port_id[3]), 
            .O(n10637));
    defparam n14717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13117 (.I0(port_id[2]), .I1(n10259), .I2(n10274), 
            .I3(port_id[3]), .O(n14717));
    defparam port_id_2__bdd_4_lut_13117.LUT_INIT = 16'he4aa;
    SB_LUT4 n14723_bdd_4_lut (.I0(n14723), .I1(ram_s_37_6), .I2(ram_s_36_6), 
            .I3(port_id[1]), .O(n9167));
    defparam n14723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13067 (.I0(port_id[0]), .I1(ram_s_38_6), 
            .I2(ram_s_39_6), .I3(port_id[1]), .O(n14723));
    defparam port_id_0__bdd_4_lut_13067.LUT_INIT = 16'he4aa;
    SB_LUT4 n14729_bdd_4_lut (.I0(n14729), .I1(ram_s_233_1), .I2(ram_s_232_1), 
            .I3(port_id[1]), .O(n10634));
    defparam n14729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13072 (.I0(port_id[0]), .I1(ram_s_234_1), 
            .I2(ram_s_235_1), .I3(port_id[1]), .O(n14729));
    defparam port_id_0__bdd_4_lut_13072.LUT_INIT = 16'he4aa;
    SB_LUT4 n14735_bdd_4_lut (.I0(n14735), .I1(ram_s_89_2), .I2(ram_s_88_2), 
            .I3(port_id[1]), .O(n8957));
    defparam n14735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13077 (.I0(port_id[0]), .I1(ram_s_90_2), 
            .I2(ram_s_91_2), .I3(port_id[1]), .O(n14735));
    defparam port_id_0__bdd_4_lut_13077.LUT_INIT = 16'he4aa;
    SB_LUT4 n14741_bdd_4_lut (.I0(n14741), .I1(ram_s_237_7), .I2(ram_s_236_7), 
            .I3(port_id[1]), .O(n10631));
    defparam n14741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13082 (.I0(port_id[0]), .I1(ram_s_238_7), 
            .I2(ram_s_239_7), .I3(port_id[1]), .O(n14741));
    defparam port_id_0__bdd_4_lut_13082.LUT_INIT = 16'he4aa;
    SB_LUT4 n14747_bdd_4_lut (.I0(n14747), .I1(ram_s_161_4), .I2(ram_s_160_4), 
            .I3(port_id[1]), .O(n9884));
    defparam n14747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13087 (.I0(port_id[0]), .I1(ram_s_162_4), 
            .I2(ram_s_163_4), .I3(port_id[1]), .O(n14747));
    defparam port_id_0__bdd_4_lut_13087.LUT_INIT = 16'he4aa;
    SB_LUT4 n14753_bdd_4_lut (.I0(n14753), .I1(ram_s_81_0), .I2(ram_s_80_0), 
            .I3(port_id[1]), .O(n8951));
    defparam n14753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13092 (.I0(port_id[0]), .I1(ram_s_82_0), 
            .I2(ram_s_83_0), .I3(port_id[1]), .O(n14753));
    defparam port_id_0__bdd_4_lut_13092.LUT_INIT = 16'he4aa;
    SB_LUT4 i1383_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_92_7), .O(n1631));   // src/ram.vhd(68[19:45])
    defparam i1383_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14759_bdd_4_lut (.I0(n14759), .I1(ram_s_81_3), .I2(ram_s_80_3), 
            .I3(port_id[1]), .O(n9161));
    defparam n14759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13097 (.I0(port_id[0]), .I1(ram_s_82_3), 
            .I2(ram_s_83_3), .I3(port_id[1]), .O(n14759));
    defparam port_id_0__bdd_4_lut_13097.LUT_INIT = 16'he4aa;
    SB_LUT4 n14765_bdd_4_lut (.I0(n14765), .I1(ram_s_177_5), .I2(ram_s_176_5), 
            .I3(port_id[1]), .O(n9491));
    defparam n14765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13107 (.I0(port_id[0]), .I1(ram_s_178_5), 
            .I2(ram_s_179_5), .I3(port_id[1]), .O(n14765));
    defparam port_id_0__bdd_4_lut_13107.LUT_INIT = 16'he4aa;
    SB_LUT4 n14777_bdd_4_lut (.I0(n14777), .I1(ram_s_157_4), .I2(ram_s_156_4), 
            .I3(port_id[1]), .O(n9881));
    defparam n14777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13122 (.I0(port_id[0]), .I1(ram_s_158_4), 
            .I2(ram_s_159_4), .I3(port_id[1]), .O(n14777));
    defparam port_id_0__bdd_4_lut_13122.LUT_INIT = 16'he4aa;
    SB_LUT4 n14789_bdd_4_lut (.I0(n14789), .I1(n13466), .I2(n14150), .I3(port_id[3]), 
            .O(n10628));
    defparam n14789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13132 (.I0(port_id[2]), .I1(n11708), .I2(n14000), 
            .I3(port_id[3]), .O(n14789));
    defparam port_id_2__bdd_4_lut_13132.LUT_INIT = 16'he4aa;
    SB_LUT4 n14795_bdd_4_lut (.I0(n14795), .I1(ram_s_101_5), .I2(ram_s_100_5), 
            .I3(port_id[1]), .O(n10286));
    defparam n14795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13127 (.I0(port_id[0]), .I1(ram_s_102_5), 
            .I2(ram_s_103_5), .I3(port_id[1]), .O(n14795));
    defparam port_id_0__bdd_4_lut_13127.LUT_INIT = 16'he4aa;
    SB_LUT4 n14801_bdd_4_lut (.I0(n14801), .I1(ram_s_173_0), .I2(ram_s_172_0), 
            .I3(port_id[1]), .O(n14804));
    defparam n14801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13137 (.I0(port_id[0]), .I1(ram_s_174_0), 
            .I2(ram_s_175_0), .I3(port_id[1]), .O(n14801));
    defparam port_id_0__bdd_4_lut_13137.LUT_INIT = 16'he4aa;
    SB_LUT4 n14807_bdd_4_lut (.I0(n14807), .I1(n13580), .I2(n13946), .I3(port_id[3]), 
            .O(n9878));
    defparam n14807_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13192 (.I0(port_id[2]), .I1(n13382), .I2(n13298), 
            .I3(port_id[3]), .O(n14807));
    defparam port_id_2__bdd_4_lut_13192.LUT_INIT = 16'he4aa;
    SB_LUT4 n14813_bdd_4_lut (.I0(n14813), .I1(ram_s_57_3), .I2(ram_s_56_3), 
            .I3(port_id[1]), .O(n8945));
    defparam n14813_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13142 (.I0(port_id[0]), .I1(ram_s_58_3), 
            .I2(ram_s_59_3), .I3(port_id[1]), .O(n14813));
    defparam port_id_0__bdd_4_lut_13142.LUT_INIT = 16'he4aa;
    SB_LUT4 n14819_bdd_4_lut (.I0(n14819), .I1(ram_s_229_1), .I2(ram_s_228_1), 
            .I3(port_id[1]), .O(n10625));
    defparam n14819_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13147 (.I0(port_id[0]), .I1(ram_s_230_1), 
            .I2(ram_s_231_1), .I3(port_id[1]), .O(n14819));
    defparam port_id_0__bdd_4_lut_13147.LUT_INIT = 16'he4aa;
    SB_LUT4 n14825_bdd_4_lut (.I0(n14825), .I1(ram_s_229_5), .I2(ram_s_228_5), 
            .I3(port_id[1]), .O(n10283));
    defparam n14825_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13152 (.I0(port_id[0]), .I1(ram_s_230_5), 
            .I2(ram_s_231_5), .I3(port_id[1]), .O(n14825));
    defparam port_id_0__bdd_4_lut_13152.LUT_INIT = 16'he4aa;
    SB_LUT4 i1382_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_92_6), .O(n1630));   // src/ram.vhd(68[19:45])
    defparam i1382_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14831_bdd_4_lut (.I0(n14831), .I1(ram_s_49_7), .I2(ram_s_48_7), 
            .I3(port_id[1]), .O(n9479));
    defparam n14831_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13157 (.I0(port_id[0]), .I1(ram_s_50_7), 
            .I2(ram_s_51_7), .I3(port_id[1]), .O(n14831));
    defparam port_id_0__bdd_4_lut_13157.LUT_INIT = 16'he4aa;
    SB_LUT4 n14837_bdd_4_lut (.I0(n14837), .I1(ram_s_225_1), .I2(ram_s_224_1), 
            .I3(port_id[1]), .O(n10622));
    defparam n14837_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13162 (.I0(port_id[0]), .I1(ram_s_226_1), 
            .I2(ram_s_227_1), .I3(port_id[1]), .O(n14837));
    defparam port_id_0__bdd_4_lut_13162.LUT_INIT = 16'he4aa;
    SB_LUT4 n14843_bdd_4_lut (.I0(n14843), .I1(ram_s_73_1), .I2(ram_s_72_1), 
            .I3(port_id[1]), .O(n10277));
    defparam n14843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13167 (.I0(port_id[0]), .I1(ram_s_74_1), 
            .I2(ram_s_75_1), .I3(port_id[1]), .O(n14843));
    defparam port_id_0__bdd_4_lut_13167.LUT_INIT = 16'he4aa;
    SB_LUT4 n14849_bdd_4_lut (.I0(n14849), .I1(ram_s_201_6), .I2(ram_s_200_6), 
            .I3(port_id[1]), .O(n9875));
    defparam n14849_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13172 (.I0(port_id[0]), .I1(ram_s_202_6), 
            .I2(ram_s_203_6), .I3(port_id[1]), .O(n14849));
    defparam port_id_0__bdd_4_lut_13172.LUT_INIT = 16'he4aa;
    SB_LUT4 n14855_bdd_4_lut (.I0(n14855), .I1(ram_s_33_6), .I2(ram_s_32_6), 
            .I3(port_id[1]), .O(n9152));
    defparam n14855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13177 (.I0(port_id[0]), .I1(ram_s_34_6), 
            .I2(ram_s_35_6), .I3(port_id[1]), .O(n14855));
    defparam port_id_0__bdd_4_lut_13177.LUT_INIT = 16'he4aa;
    SB_LUT4 n14861_bdd_4_lut (.I0(n14861), .I1(ram_s_221_3), .I2(ram_s_220_3), 
            .I3(port_id[1]), .O(n10274));
    defparam n14861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13182 (.I0(port_id[0]), .I1(ram_s_222_3), 
            .I2(ram_s_223_3), .I3(port_id[1]), .O(n14861));
    defparam port_id_0__bdd_4_lut_13182.LUT_INIT = 16'he4aa;
    SB_LUT4 n14867_bdd_4_lut (.I0(n14867), .I1(ram_s_153_4), .I2(ram_s_152_4), 
            .I3(port_id[1]), .O(n9872));
    defparam n14867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13187 (.I0(port_id[0]), .I1(ram_s_154_4), 
            .I2(ram_s_155_4), .I3(port_id[1]), .O(n14867));
    defparam port_id_0__bdd_4_lut_13187.LUT_INIT = 16'he4aa;
    SB_LUT4 n14873_bdd_4_lut (.I0(n14873), .I1(ram_s_69_1), .I2(ram_s_68_1), 
            .I3(port_id[1]), .O(n10271));
    defparam n14873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13197 (.I0(port_id[0]), .I1(ram_s_70_1), 
            .I2(ram_s_71_1), .I3(port_id[1]), .O(n14873));
    defparam port_id_0__bdd_4_lut_13197.LUT_INIT = 16'he4aa;
    SB_LUT4 n14879_bdd_4_lut (.I0(n14879), .I1(n9824), .I2(n9812), .I3(port_id[3]), 
            .O(n10268));
    defparam n14879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13207 (.I0(port_id[2]), .I1(n9830), .I2(n9851), 
            .I3(port_id[3]), .O(n14879));
    defparam port_id_2__bdd_4_lut_13207.LUT_INIT = 16'he4aa;
    SB_LUT4 n14885_bdd_4_lut (.I0(n14885), .I1(ram_s_121_5), .I2(ram_s_120_5), 
            .I3(port_id[1]), .O(n10619));
    defparam n14885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13202 (.I0(port_id[0]), .I1(ram_s_122_5), 
            .I2(ram_s_123_5), .I3(port_id[1]), .O(n14885));
    defparam port_id_0__bdd_4_lut_13202.LUT_INIT = 16'he4aa;
    SB_LUT4 n14891_bdd_4_lut (.I0(n14891), .I1(ram_s_161_3), .I2(ram_s_160_3), 
            .I3(port_id[1]), .O(n14894));
    defparam n14891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13217 (.I0(port_id[0]), .I1(ram_s_162_3), 
            .I2(ram_s_163_3), .I3(port_id[1]), .O(n14891));
    defparam port_id_0__bdd_4_lut_13217.LUT_INIT = 16'he4aa;
    SB_LUT4 n14897_bdd_4_lut (.I0(n14897), .I1(n12284), .I2(n12398), .I3(port_id[3]), 
            .O(n10616));
    defparam n14897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13277 (.I0(port_id[2]), .I1(n12008), .I2(n11612), 
            .I3(port_id[3]), .O(n14897));
    defparam port_id_2__bdd_4_lut_13277.LUT_INIT = 16'he4aa;
    SB_LUT4 i1381_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_92_5), .O(n1629));   // src/ram.vhd(68[19:45])
    defparam i1381_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14909_bdd_4_lut (.I0(n14909), .I1(ram_s_149_4), .I2(ram_s_148_4), 
            .I3(port_id[1]), .O(n9863));
    defparam n14909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13222 (.I0(port_id[0]), .I1(ram_s_150_4), 
            .I2(ram_s_151_4), .I3(port_id[1]), .O(n14909));
    defparam port_id_0__bdd_4_lut_13222.LUT_INIT = 16'he4aa;
    SB_LUT4 n14915_bdd_4_lut (.I0(n14915), .I1(ram_s_197_6), .I2(ram_s_196_6), 
            .I3(port_id[1]), .O(n9860));
    defparam n14915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13227 (.I0(port_id[0]), .I1(ram_s_198_6), 
            .I2(ram_s_199_6), .I3(port_id[1]), .O(n14915));
    defparam port_id_0__bdd_4_lut_13227.LUT_INIT = 16'he4aa;
    SB_LUT4 n14921_bdd_4_lut (.I0(n14921), .I1(ram_s_233_7), .I2(ram_s_232_7), 
            .I3(port_id[1]), .O(n10613));
    defparam n14921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13232 (.I0(port_id[0]), .I1(ram_s_234_7), 
            .I2(ram_s_235_7), .I3(port_id[1]), .O(n14921));
    defparam port_id_0__bdd_4_lut_13232.LUT_INIT = 16'he4aa;
    SB_LUT4 n14927_bdd_4_lut (.I0(n14927), .I1(ram_s_169_0), .I2(ram_s_168_0), 
            .I3(port_id[1]), .O(n14930));
    defparam n14927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13242 (.I0(port_id[0]), .I1(ram_s_170_0), 
            .I2(ram_s_171_0), .I3(port_id[1]), .O(n14927));
    defparam port_id_0__bdd_4_lut_13242.LUT_INIT = 16'he4aa;
    SB_LUT4 n14933_bdd_4_lut (.I0(n14933), .I1(n11690), .I2(n8843), .I3(port_id[7]), 
            .O(spm_ram_data[4]));
    defparam n14933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_6__bdd_4_lut (.I0(port_id[6]), .I1(n11528), .I2(n11174), 
            .I3(port_id[7]), .O(n14933));
    defparam port_id_6__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14939_bdd_4_lut (.I0(n14939), .I1(ram_s_77_0), .I2(ram_s_76_0), 
            .I3(port_id[1]), .O(n8939));
    defparam n14939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13247 (.I0(port_id[0]), .I1(ram_s_78_0), 
            .I2(ram_s_79_0), .I3(port_id[1]), .O(n14939));
    defparam port_id_0__bdd_4_lut_13247.LUT_INIT = 16'he4aa;
    SB_LUT4 n14945_bdd_4_lut (.I0(n14945), .I1(ram_s_217_3), .I2(ram_s_216_3), 
            .I3(port_id[1]), .O(n10259));
    defparam n14945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13252 (.I0(port_id[0]), .I1(ram_s_218_3), 
            .I2(ram_s_219_3), .I3(port_id[1]), .O(n14945));
    defparam port_id_0__bdd_4_lut_13252.LUT_INIT = 16'he4aa;
    SB_LUT4 n14951_bdd_4_lut (.I0(n14951), .I1(ram_s_25_5), .I2(ram_s_24_5), 
            .I3(port_id[1]), .O(n9467));
    defparam n14951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13257 (.I0(port_id[0]), .I1(ram_s_26_5), 
            .I2(ram_s_27_5), .I3(port_id[1]), .O(n14951));
    defparam port_id_0__bdd_4_lut_13257.LUT_INIT = 16'he4aa;
    SB_LUT4 n14957_bdd_4_lut (.I0(n14957), .I1(ram_s_221_1), .I2(ram_s_220_1), 
            .I3(port_id[1]), .O(n10610));
    defparam n14957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13262 (.I0(port_id[0]), .I1(ram_s_222_1), 
            .I2(ram_s_223_1), .I3(port_id[1]), .O(n14957));
    defparam port_id_0__bdd_4_lut_13262.LUT_INIT = 16'he4aa;
    SB_LUT4 n14963_bdd_4_lut (.I0(n14963), .I1(ram_s_65_5), .I2(ram_s_64_5), 
            .I3(port_id[1]), .O(n9140));
    defparam n14963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13272 (.I0(port_id[0]), .I1(ram_s_66_5), 
            .I2(ram_s_67_5), .I3(port_id[1]), .O(n14963));
    defparam port_id_0__bdd_4_lut_13272.LUT_INIT = 16'he4aa;
    SB_LUT4 n14975_bdd_4_lut (.I0(n14975), .I1(ram_s_145_4), .I2(ram_s_144_4), 
            .I3(port_id[1]), .O(n9854));
    defparam n14975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13282 (.I0(port_id[0]), .I1(ram_s_146_4), 
            .I2(ram_s_147_4), .I3(port_id[1]), .O(n14975));
    defparam port_id_0__bdd_4_lut_13282.LUT_INIT = 16'he4aa;
    SB_LUT4 n14981_bdd_4_lut (.I0(n14981), .I1(n13550), .I2(n13760), .I3(port_id[3]), 
            .O(n10607));
    defparam n14981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13322 (.I0(port_id[2]), .I1(n12968), .I2(n12716), 
            .I3(port_id[3]), .O(n14981));
    defparam port_id_2__bdd_4_lut_13322.LUT_INIT = 16'he4aa;
    SB_LUT4 n14987_bdd_4_lut (.I0(n14987), .I1(ram_s_65_1), .I2(ram_s_64_1), 
            .I3(port_id[1]), .O(n10256));
    defparam n14987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13287 (.I0(port_id[0]), .I1(ram_s_66_1), 
            .I2(ram_s_67_1), .I3(port_id[1]), .O(n14987));
    defparam port_id_0__bdd_4_lut_13287.LUT_INIT = 16'he4aa;
    SB_LUT4 n14993_bdd_4_lut (.I0(n14993), .I1(ram_s_117_3), .I2(ram_s_116_3), 
            .I3(port_id[1]), .O(n9461));
    defparam n14993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13292 (.I0(port_id[0]), .I1(ram_s_118_3), 
            .I2(ram_s_119_3), .I3(port_id[1]), .O(n14993));
    defparam port_id_0__bdd_4_lut_13292.LUT_INIT = 16'he4aa;
    SB_LUT4 n14999_bdd_4_lut (.I0(n14999), .I1(ram_s_205_2), .I2(ram_s_204_2), 
            .I3(port_id[1]), .O(n9458));
    defparam n14999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13297 (.I0(port_id[0]), .I1(ram_s_206_2), 
            .I2(ram_s_207_2), .I3(port_id[1]), .O(n14999));
    defparam port_id_0__bdd_4_lut_13297.LUT_INIT = 16'he4aa;
    SB_LUT4 n15005_bdd_4_lut (.I0(n15005), .I1(ram_s_141_4), .I2(ram_s_140_4), 
            .I3(port_id[1]), .O(n9851));
    defparam n15005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13302 (.I0(port_id[0]), .I1(ram_s_142_4), 
            .I2(ram_s_143_4), .I3(port_id[1]), .O(n15005));
    defparam port_id_0__bdd_4_lut_13302.LUT_INIT = 16'he4aa;
    SB_LUT4 n15011_bdd_4_lut (.I0(n15011), .I1(ram_s_217_1), .I2(ram_s_216_1), 
            .I3(port_id[1]), .O(n10604));
    defparam n15011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13307 (.I0(port_id[0]), .I1(ram_s_218_1), 
            .I2(ram_s_219_1), .I3(port_id[1]), .O(n15011));
    defparam port_id_0__bdd_4_lut_13307.LUT_INIT = 16'he4aa;
    SB_LUT4 n15017_bdd_4_lut (.I0(n15017), .I1(ram_s_61_1), .I2(ram_s_60_1), 
            .I3(port_id[1]), .O(n10253));
    defparam n15017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13317 (.I0(port_id[0]), .I1(ram_s_62_1), 
            .I2(ram_s_63_1), .I3(port_id[1]), .O(n15017));
    defparam port_id_0__bdd_4_lut_13317.LUT_INIT = 16'he4aa;
    SB_LUT4 n15029_bdd_4_lut (.I0(n15029), .I1(ram_s_85_5), .I2(ram_s_84_5), 
            .I3(port_id[1]), .O(n9842));
    defparam n15029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13327 (.I0(port_id[0]), .I1(ram_s_86_5), 
            .I2(ram_s_87_5), .I3(port_id[1]), .O(n15029));
    defparam port_id_0__bdd_4_lut_13327.LUT_INIT = 16'he4aa;
    SB_LUT4 n15035_bdd_4_lut (.I0(n15035), .I1(n13454), .I2(n13640), .I3(port_id[3]), 
            .O(n10250));
    defparam n15035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13357 (.I0(port_id[2]), .I1(n13376), .I2(n13214), 
            .I3(port_id[3]), .O(n15035));
    defparam port_id_2__bdd_4_lut_13357.LUT_INIT = 16'he4aa;
    SB_LUT4 n15041_bdd_4_lut (.I0(n15041), .I1(ram_s_229_7), .I2(ram_s_228_7), 
            .I3(port_id[1]), .O(n10601));
    defparam n15041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13332 (.I0(port_id[0]), .I1(ram_s_230_7), 
            .I2(ram_s_231_7), .I3(port_id[1]), .O(n15041));
    defparam port_id_0__bdd_4_lut_13332.LUT_INIT = 16'he4aa;
    SB_LUT4 n15047_bdd_4_lut (.I0(n15047), .I1(ram_s_201_2), .I2(ram_s_200_2), 
            .I3(port_id[1]), .O(n9449));
    defparam n15047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13337 (.I0(port_id[0]), .I1(ram_s_202_2), 
            .I2(ram_s_203_2), .I3(port_id[1]), .O(n15047));
    defparam port_id_0__bdd_4_lut_13337.LUT_INIT = 16'he4aa;
    SB_LUT4 n15053_bdd_4_lut (.I0(n15053), .I1(ram_s_29_6), .I2(ram_s_28_6), 
            .I3(port_id[1]), .O(n9131));
    defparam n15053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13342 (.I0(port_id[0]), .I1(ram_s_30_6), 
            .I2(ram_s_31_6), .I3(port_id[1]), .O(n15053));
    defparam port_id_0__bdd_4_lut_13342.LUT_INIT = 16'he4aa;
    SB_LUT4 n15059_bdd_4_lut (.I0(n15059), .I1(ram_s_197_5), .I2(ram_s_196_5), 
            .I3(port_id[1]), .O(n15062));
    defparam n15059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13347 (.I0(port_id[0]), .I1(ram_s_198_5), 
            .I2(ram_s_199_5), .I3(port_id[1]), .O(n15059));
    defparam port_id_0__bdd_4_lut_13347.LUT_INIT = 16'he4aa;
    SB_LUT4 n15065_bdd_4_lut (.I0(n15065), .I1(ram_s_225_5), .I2(ram_s_224_5), 
            .I3(port_id[1]), .O(n10247));
    defparam n15065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13352 (.I0(port_id[0]), .I1(ram_s_226_5), 
            .I2(ram_s_227_5), .I3(port_id[1]), .O(n15065));
    defparam port_id_0__bdd_4_lut_13352.LUT_INIT = 16'he4aa;
    SB_LUT4 n15071_bdd_4_lut (.I0(n15071), .I1(ram_s_85_2), .I2(ram_s_84_2), 
            .I3(port_id[1]), .O(n8933));
    defparam n15071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13362 (.I0(port_id[0]), .I1(ram_s_86_2), 
            .I2(ram_s_87_2), .I3(port_id[1]), .O(n15071));
    defparam port_id_0__bdd_4_lut_13362.LUT_INIT = 16'he4aa;
    SB_LUT4 n15077_bdd_4_lut (.I0(n15077), .I1(n14432), .I2(n14624), .I3(port_id[3]), 
            .O(n10598));
    defparam n15077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13412 (.I0(port_id[2]), .I1(n14288), .I2(n14102), 
            .I3(port_id[3]), .O(n15077));
    defparam port_id_2__bdd_4_lut_13412.LUT_INIT = 16'he4aa;
    SB_LUT4 n15083_bdd_4_lut (.I0(n15083), .I1(ram_s_73_0), .I2(ram_s_72_0), 
            .I3(port_id[1]), .O(n8930));
    defparam n15083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13367 (.I0(port_id[0]), .I1(ram_s_74_0), 
            .I2(ram_s_75_0), .I3(port_id[1]), .O(n15083));
    defparam port_id_0__bdd_4_lut_13367.LUT_INIT = 16'he4aa;
    SB_LUT4 n15089_bdd_4_lut (.I0(n15089), .I1(ram_s_157_0), .I2(ram_s_156_0), 
            .I3(port_id[1]), .O(n9122));
    defparam n15089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13372 (.I0(port_id[0]), .I1(ram_s_158_0), 
            .I2(ram_s_159_0), .I3(port_id[1]), .O(n15089));
    defparam port_id_0__bdd_4_lut_13372.LUT_INIT = 16'he4aa;
    SB_LUT4 i1380_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_92_4), .O(n1628));   // src/ram.vhd(68[19:45])
    defparam i1380_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15095_bdd_4_lut (.I0(n15095), .I1(ram_s_113_3), .I2(ram_s_112_3), 
            .I3(port_id[1]), .O(n9440));
    defparam n15095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13377 (.I0(port_id[0]), .I1(ram_s_114_3), 
            .I2(ram_s_115_3), .I3(port_id[1]), .O(n15095));
    defparam port_id_0__bdd_4_lut_13377.LUT_INIT = 16'he4aa;
    SB_LUT4 n15101_bdd_4_lut (.I0(n15101), .I1(ram_s_5_3), .I2(ram_s_4_3), 
            .I3(port_id[1]), .O(n10595));
    defparam n15101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13382 (.I0(port_id[0]), .I1(ram_s_6_3), 
            .I2(ram_s_7_3), .I3(port_id[1]), .O(n15101));
    defparam port_id_0__bdd_4_lut_13382.LUT_INIT = 16'he4aa;
    SB_LUT4 n15107_bdd_4_lut (.I0(n15107), .I1(ram_s_193_6), .I2(ram_s_192_6), 
            .I3(port_id[1]), .O(n9833));
    defparam n15107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13387 (.I0(port_id[0]), .I1(ram_s_194_6), 
            .I2(ram_s_195_6), .I3(port_id[1]), .O(n15107));
    defparam port_id_0__bdd_4_lut_13387.LUT_INIT = 16'he4aa;
    SB_LUT4 n15113_bdd_4_lut (.I0(n15113), .I1(ram_s_25_6), .I2(ram_s_24_6), 
            .I3(port_id[1]), .O(n9119));
    defparam n15113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13392 (.I0(port_id[0]), .I1(ram_s_26_6), 
            .I2(ram_s_27_6), .I3(port_id[1]), .O(n15113));
    defparam port_id_0__bdd_4_lut_13392.LUT_INIT = 16'he4aa;
    SB_LUT4 n15119_bdd_4_lut (.I0(n15119), .I1(ram_s_137_4), .I2(ram_s_136_4), 
            .I3(port_id[1]), .O(n9830));
    defparam n15119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13397 (.I0(port_id[0]), .I1(ram_s_138_4), 
            .I2(ram_s_139_4), .I3(port_id[1]), .O(n15119));
    defparam port_id_0__bdd_4_lut_13397.LUT_INIT = 16'he4aa;
    SB_LUT4 n15125_bdd_4_lut (.I0(n15125), .I1(ram_s_149_7), .I2(ram_s_148_7), 
            .I3(port_id[1]), .O(n15128));
    defparam n15125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13402 (.I0(port_id[0]), .I1(ram_s_150_7), 
            .I2(ram_s_151_7), .I3(port_id[1]), .O(n15125));
    defparam port_id_0__bdd_4_lut_13402.LUT_INIT = 16'he4aa;
    SB_LUT4 n15131_bdd_4_lut (.I0(n15131), .I1(ram_s_77_3), .I2(ram_s_76_3), 
            .I3(port_id[1]), .O(n9116));
    defparam n15131_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13407 (.I0(port_id[0]), .I1(ram_s_78_3), 
            .I2(ram_s_79_3), .I3(port_id[1]), .O(n15131));
    defparam port_id_0__bdd_4_lut_13407.LUT_INIT = 16'he4aa;
    SB_LUT4 n15137_bdd_4_lut (.I0(n15137), .I1(ram_s_45_7), .I2(ram_s_44_7), 
            .I3(port_id[1]), .O(n9437));
    defparam n15137_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13417 (.I0(port_id[0]), .I1(ram_s_46_7), 
            .I2(ram_s_47_7), .I3(port_id[1]), .O(n15137));
    defparam port_id_0__bdd_4_lut_13417.LUT_INIT = 16'he4aa;
    SB_LUT4 n15143_bdd_4_lut (.I0(n15143), .I1(n12800), .I2(n13022), .I3(port_id[3]), 
            .O(n9827));
    defparam n15143_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13427 (.I0(port_id[2]), .I1(n9104), .I2(n9113), 
            .I3(port_id[3]), .O(n15143));
    defparam port_id_2__bdd_4_lut_13427.LUT_INIT = 16'he4aa;
    SB_LUT4 n15149_bdd_4_lut (.I0(n15149), .I1(ram_s_57_1), .I2(ram_s_56_1), 
            .I3(port_id[1]), .O(n10241));
    defparam n15149_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13422 (.I0(port_id[0]), .I1(ram_s_58_1), 
            .I2(ram_s_59_1), .I3(port_id[1]), .O(n15149));
    defparam port_id_0__bdd_4_lut_13422.LUT_INIT = 16'he4aa;
    SB_LUT4 n15155_bdd_4_lut (.I0(n15155), .I1(ram_s_69_0), .I2(ram_s_68_0), 
            .I3(port_id[1]), .O(n8927));
    defparam n15155_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13432 (.I0(port_id[0]), .I1(ram_s_70_0), 
            .I2(ram_s_71_0), .I3(port_id[1]), .O(n15155));
    defparam port_id_0__bdd_4_lut_13432.LUT_INIT = 16'he4aa;
    SB_LUT4 n15161_bdd_4_lut (.I0(n15161), .I1(n10238), .I2(n12464), .I3(port_id[3]), 
            .O(n10592));
    defparam n15161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13462 (.I0(port_id[2]), .I1(n11624), .I2(n12050), 
            .I3(port_id[3]), .O(n15161));
    defparam port_id_2__bdd_4_lut_13462.LUT_INIT = 16'he4aa;
    SB_LUT4 i1379_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_92_3), .O(n1627));   // src/ram.vhd(68[19:45])
    defparam i1379_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n15167_bdd_4_lut (.I0(n15167), .I1(ram_s_125_2), .I2(ram_s_124_2), 
            .I3(port_id[1]), .O(n9113));
    defparam n15167_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13437 (.I0(port_id[0]), .I1(ram_s_126_2), 
            .I2(ram_s_127_2), .I3(port_id[1]), .O(n15167));
    defparam port_id_0__bdd_4_lut_13437.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i159_2_lut (.I0(n96_adj_864), .I1(port_id[6]), 
            .I2(wea[0]), .I3(wea[0]), .O(n159));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n15173_bdd_4_lut (.I0(n15173), .I1(ram_s_133_4), .I2(ram_s_132_4), 
            .I3(port_id[1]), .O(n9824));
    defparam n15173_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13442 (.I0(port_id[0]), .I1(ram_s_134_4), 
            .I2(ram_s_135_4), .I3(port_id[1]), .O(n15173));
    defparam port_id_0__bdd_4_lut_13442.LUT_INIT = 16'he4aa;
    SB_LUT4 n15179_bdd_4_lut (.I0(n15179), .I1(ram_s_213_1), .I2(ram_s_212_1), 
            .I3(port_id[1]), .O(n10589));
    defparam n15179_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13447 (.I0(port_id[0]), .I1(ram_s_214_1), 
            .I2(ram_s_215_1), .I3(port_id[1]), .O(n15179));
    defparam port_id_0__bdd_4_lut_13447.LUT_INIT = 16'he4aa;
    SB_LUT4 n15185_bdd_4_lut (.I0(n15185), .I1(ram_s_153_0), .I2(ram_s_152_0), 
            .I3(port_id[1]), .O(n9110));
    defparam n15185_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13452 (.I0(port_id[0]), .I1(ram_s_154_0), 
            .I2(ram_s_155_0), .I3(port_id[1]), .O(n15185));
    defparam port_id_0__bdd_4_lut_13452.LUT_INIT = 16'he4aa;
    SB_LUT4 n15191_bdd_4_lut (.I0(n15191), .I1(ram_s_149_0), .I2(ram_s_148_0), 
            .I3(port_id[1]), .O(n9107));
    defparam n15191_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13457 (.I0(port_id[0]), .I1(ram_s_150_0), 
            .I2(ram_s_151_0), .I3(port_id[1]), .O(n15191));
    defparam port_id_0__bdd_4_lut_13457.LUT_INIT = 16'he4aa;
    SB_LUT4 n15197_bdd_4_lut (.I0(n15197), .I1(ram_s_209_1), .I2(ram_s_208_1), 
            .I3(port_id[1]), .O(n10586));
    defparam n15197_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13467 (.I0(port_id[0]), .I1(ram_s_210_1), 
            .I2(ram_s_211_1), .I3(port_id[1]), .O(n15197));
    defparam port_id_0__bdd_4_lut_13467.LUT_INIT = 16'he4aa;
    SB_LUT4 n15203_bdd_4_lut (.I0(n15203), .I1(n14702), .I2(n14894), .I3(port_id[3]), 
            .O(n10583));
    defparam n15203_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut_13522 (.I0(port_id[2]), .I1(n14384), .I2(n14126), 
            .I3(port_id[3]), .O(n15203));
    defparam port_id_2__bdd_4_lut_13522.LUT_INIT = 16'he4aa;
    SB_LUT4 n15209_bdd_4_lut (.I0(n15209), .I1(ram_s_145_5), .I2(ram_s_144_5), 
            .I3(port_id[1]), .O(n15212));
    defparam n15209_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13472 (.I0(port_id[0]), .I1(ram_s_146_5), 
            .I2(ram_s_147_5), .I3(port_id[1]), .O(n15209));
    defparam port_id_0__bdd_4_lut_13472.LUT_INIT = 16'he4aa;
    SB_LUT4 n15215_bdd_4_lut (.I0(n15215), .I1(ram_s_81_2), .I2(ram_s_80_2), 
            .I3(port_id[1]), .O(n8921));
    defparam n15215_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13477 (.I0(port_id[0]), .I1(ram_s_82_2), 
            .I2(ram_s_83_2), .I3(port_id[1]), .O(n15215));
    defparam port_id_0__bdd_4_lut_13477.LUT_INIT = 16'he4aa;
    SB_LUT4 n15221_bdd_4_lut (.I0(n15221), .I1(ram_s_37_5), .I2(ram_s_36_5), 
            .I3(port_id[1]), .O(n10238));
    defparam n15221_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13482 (.I0(port_id[0]), .I1(ram_s_38_5), 
            .I2(ram_s_39_5), .I3(port_id[1]), .O(n15221));
    defparam port_id_0__bdd_4_lut_13482.LUT_INIT = 16'he4aa;
    SB_LUT4 n15227_bdd_4_lut (.I0(n15227), .I1(ram_s_189_6), .I2(ram_s_188_6), 
            .I3(port_id[1]), .O(n9821));
    defparam n15227_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13487 (.I0(port_id[0]), .I1(ram_s_190_6), 
            .I2(ram_s_191_6), .I3(port_id[1]), .O(n15227));
    defparam port_id_0__bdd_4_lut_13487.LUT_INIT = 16'he4aa;
    SB_LUT4 n15233_bdd_4_lut (.I0(n15233), .I1(ram_s_225_7), .I2(ram_s_224_7), 
            .I3(port_id[1]), .O(n10580));
    defparam n15233_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13497 (.I0(port_id[0]), .I1(ram_s_226_7), 
            .I2(ram_s_227_7), .I3(port_id[1]), .O(n15233));
    defparam port_id_0__bdd_4_lut_13497.LUT_INIT = 16'he4aa;
    SB_LUT4 i1378_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_92_2), .O(n1626));   // src/ram.vhd(68[19:45])
    defparam i1378_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i161_2_lut (.I0(n98), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n161));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n15245_bdd_4_lut (.I0(n15245), .I1(ram_s_157_3), .I2(ram_s_156_3), 
            .I3(port_id[1]), .O(n9818));
    defparam n15245_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13502 (.I0(port_id[0]), .I1(ram_s_158_3), 
            .I2(ram_s_159_3), .I3(port_id[1]), .O(n15245));
    defparam port_id_0__bdd_4_lut_13502.LUT_INIT = 16'he4aa;
    SB_LUT4 n15251_bdd_4_lut (.I0(n15251), .I1(ram_s_205_1), .I2(ram_s_204_1), 
            .I3(port_id[1]), .O(n10577));
    defparam n15251_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13507 (.I0(port_id[0]), .I1(ram_s_206_1), 
            .I2(ram_s_207_1), .I3(port_id[1]), .O(n15251));
    defparam port_id_0__bdd_4_lut_13507.LUT_INIT = 16'he4aa;
    SB_LUT4 n15257_bdd_4_lut (.I0(n15257), .I1(ram_s_213_3), .I2(ram_s_212_3), 
            .I3(port_id[1]), .O(n10232));
    defparam n15257_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13512 (.I0(port_id[0]), .I1(ram_s_214_3), 
            .I2(ram_s_215_3), .I3(port_id[1]), .O(n15257));
    defparam port_id_0__bdd_4_lut_13512.LUT_INIT = 16'he4aa;
    SB_LUT4 n15263_bdd_4_lut (.I0(n15263), .I1(ram_s_129_4), .I2(ram_s_128_4), 
            .I3(port_id[1]), .O(n9812));
    defparam n15263_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13517 (.I0(port_id[0]), .I1(ram_s_130_4), 
            .I2(ram_s_131_4), .I3(port_id[1]), .O(n15263));
    defparam port_id_0__bdd_4_lut_13517.LUT_INIT = 16'he4aa;
    SB_LUT4 n15269_bdd_4_lut (.I0(n15269), .I1(ram_s_125_4), .I2(ram_s_124_4), 
            .I3(port_id[1]), .O(n9809));
    defparam n15269_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13527 (.I0(port_id[0]), .I1(ram_s_126_4), 
            .I2(ram_s_127_4), .I3(port_id[1]), .O(n15269));
    defparam port_id_0__bdd_4_lut_13527.LUT_INIT = 16'he4aa;
    SB_LUT4 n15275_bdd_4_lut (.I0(n15275), .I1(n13610), .I2(n14084), .I3(port_id[3]), 
            .O(n9806));
    defparam n15275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_2__bdd_4_lut (.I0(port_id[2]), .I1(n13346), .I2(n13250), 
            .I3(port_id[3]), .O(n15275));
    defparam port_id_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n15281_bdd_4_lut (.I0(n15281), .I1(ram_s_197_2), .I2(ram_s_196_2), 
            .I3(port_id[1]), .O(n9428));
    defparam n15281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13532 (.I0(port_id[0]), .I1(ram_s_198_2), 
            .I2(ram_s_199_2), .I3(port_id[1]), .O(n15281));
    defparam port_id_0__bdd_4_lut_13532.LUT_INIT = 16'he4aa;
    SB_LUT4 n15287_bdd_4_lut (.I0(n15287), .I1(ram_s_121_2), .I2(ram_s_120_2), 
            .I3(port_id[1]), .O(n9104));
    defparam n15287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13537 (.I0(port_id[0]), .I1(ram_s_122_2), 
            .I2(ram_s_123_2), .I3(port_id[1]), .O(n15287));
    defparam port_id_0__bdd_4_lut_13537.LUT_INIT = 16'he4aa;
    SB_LUT4 n15293_bdd_4_lut (.I0(n15293), .I1(ram_s_185_6), .I2(ram_s_184_6), 
            .I3(port_id[1]), .O(n9803));
    defparam n15293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13542 (.I0(port_id[0]), .I1(ram_s_186_6), 
            .I2(ram_s_187_6), .I3(port_id[1]), .O(n15293));
    defparam port_id_0__bdd_4_lut_13542.LUT_INIT = 16'he4aa;
    SB_LUT4 n15299_bdd_4_lut (.I0(n15299), .I1(ram_s_21_6), .I2(ram_s_20_6), 
            .I3(port_id[1]), .O(n9101));
    defparam n15299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13547 (.I0(port_id[0]), .I1(ram_s_22_6), 
            .I2(ram_s_23_6), .I3(port_id[1]), .O(n15299));
    defparam port_id_0__bdd_4_lut_13547.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i163_2_lut (.I0(n100), .I1(port_id[6]), .I2(wea[0]), 
            .I3(wea[0]), .O(n163));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n15305_bdd_4_lut (.I0(n15305), .I1(ram_s_53_1), .I2(ram_s_52_1), 
            .I3(port_id[1]), .O(n10229));
    defparam n15305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13552 (.I0(port_id[0]), .I1(ram_s_54_1), 
            .I2(ram_s_55_1), .I3(port_id[1]), .O(n15305));
    defparam port_id_0__bdd_4_lut_13552.LUT_INIT = 16'he4aa;
    SB_LUT4 n15311_bdd_4_lut (.I0(n15311), .I1(ram_s_1_3), .I2(ram_s_0_3), 
            .I3(port_id[1]), .O(n10574));
    defparam n15311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut_13557 (.I0(port_id[0]), .I1(ram_s_2_3), 
            .I2(ram_s_3_3), .I3(port_id[1]), .O(n15311));
    defparam port_id_0__bdd_4_lut_13557.LUT_INIT = 16'he4aa;
    SB_LUT4 n15317_bdd_4_lut (.I0(n15317), .I1(ram_s_145_0), .I2(ram_s_144_0), 
            .I3(port_id[1]), .O(n9098));
    defparam n15317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_0__bdd_4_lut (.I0(port_id[0]), .I1(ram_s_146_0), .I2(ram_s_147_0), 
            .I3(port_id[1]), .O(n15317));
    defparam port_id_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1377_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_92_1), .O(n1625));   // src/ram.vhd(68[19:45])
    defparam i1377_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1376_3_lut_4_lut (.I0(n191_adj_861), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_92_0), .O(n1624));   // src/ram.vhd(68[19:45])
    defparam i1376_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i180_2_lut_3_lut (.I0(n51), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n180));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i180_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i179_2_lut_3_lut (.I0(n51), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n179));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i179_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1375_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_91_7), .O(n1623));   // src/ram.vhd(68[19:45])
    defparam i1375_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1374_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_91_6), .O(n1622));   // src/ram.vhd(68[19:45])
    defparam i1374_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1373_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_91_5), .O(n1621));   // src/ram.vhd(68[19:45])
    defparam i1373_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1372_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_91_4), .O(n1620));   // src/ram.vhd(68[19:45])
    defparam i1372_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1371_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_91_3), .O(n1619));   // src/ram.vhd(68[19:45])
    defparam i1371_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1370_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_91_2), .O(n1618));   // src/ram.vhd(68[19:45])
    defparam i1370_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1369_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_91_1), .O(n1617));   // src/ram.vhd(68[19:45])
    defparam i1369_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1368_3_lut_4_lut (.I0(n189_adj_882), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_91_0), .O(n1616));   // src/ram.vhd(68[19:45])
    defparam i1368_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1367_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_90_7), .O(n1615));   // src/ram.vhd(68[19:45])
    defparam i1367_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1366_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_90_6), .O(n1614));   // src/ram.vhd(68[19:45])
    defparam i1366_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1365_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_90_5), .O(n1613));   // src/ram.vhd(68[19:45])
    defparam i1365_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1364_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_90_4), .O(n1612));   // src/ram.vhd(68[19:45])
    defparam i1364_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1363_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_90_3), .O(n1611));   // src/ram.vhd(68[19:45])
    defparam i1363_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1362_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_90_2), .O(n1610));   // src/ram.vhd(68[19:45])
    defparam i1362_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1361_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_90_1), .O(n1609));   // src/ram.vhd(68[19:45])
    defparam i1361_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1360_3_lut_4_lut (.I0(n187_adj_877), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_90_0), .O(n1608));   // src/ram.vhd(68[19:45])
    defparam i1360_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2351_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_213_7), .O(n2599));   // src/ram.vhd(68[19:45])
    defparam i2351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2350_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_213_6), .O(n2598));   // src/ram.vhd(68[19:45])
    defparam i2350_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2349_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_213_5), .O(n2597));   // src/ram.vhd(68[19:45])
    defparam i2349_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2348_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_213_4), .O(n2596));   // src/ram.vhd(68[19:45])
    defparam i2348_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2347_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_213_3), .O(n2595));   // src/ram.vhd(68[19:45])
    defparam i2347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2346_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_213_2), .O(n2594));   // src/ram.vhd(68[19:45])
    defparam i2346_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2345_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_213_1), .O(n2593));   // src/ram.vhd(68[19:45])
    defparam i2345_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2344_3_lut_4_lut (.I0(n177), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_213_0), .O(n2592));   // src/ram.vhd(68[19:45])
    defparam i2344_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1359_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_89_7), .O(n1607));   // src/ram.vhd(68[19:45])
    defparam i1359_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1358_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_89_6), .O(n1606));   // src/ram.vhd(68[19:45])
    defparam i1358_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1357_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_89_5), .O(n1605));   // src/ram.vhd(68[19:45])
    defparam i1357_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1356_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_89_4), .O(n1604));   // src/ram.vhd(68[19:45])
    defparam i1356_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1355_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_89_3), .O(n1603));   // src/ram.vhd(68[19:45])
    defparam i1355_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1354_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_89_2), .O(n1602));   // src/ram.vhd(68[19:45])
    defparam i1354_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1353_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_89_1), .O(n1601));   // src/ram.vhd(68[19:45])
    defparam i1353_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1352_3_lut_4_lut (.I0(n185_adj_878), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_89_0), .O(n1600));   // src/ram.vhd(68[19:45])
    defparam i1352_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1351_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_88_7), .O(n1599));   // src/ram.vhd(68[19:45])
    defparam i1351_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1350_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_88_6), .O(n1598));   // src/ram.vhd(68[19:45])
    defparam i1350_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1349_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_88_5), .O(n1597));   // src/ram.vhd(68[19:45])
    defparam i1349_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1348_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_88_4), .O(n1596));   // src/ram.vhd(68[19:45])
    defparam i1348_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1347_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_88_3), .O(n1595));   // src/ram.vhd(68[19:45])
    defparam i1347_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1346_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_88_2), .O(n1594));   // src/ram.vhd(68[19:45])
    defparam i1346_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1345_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_88_1), .O(n1593));   // src/ram.vhd(68[19:45])
    defparam i1345_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1344_3_lut_4_lut (.I0(n183_adj_883), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_88_0), .O(n1592));   // src/ram.vhd(68[19:45])
    defparam i1344_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2343_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_212_7), .O(n2591));   // src/ram.vhd(68[19:45])
    defparam i2343_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2342_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_212_6), .O(n2590));   // src/ram.vhd(68[19:45])
    defparam i2342_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2341_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_212_5), .O(n2589));   // src/ram.vhd(68[19:45])
    defparam i2341_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2340_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_212_4), .O(n2588));   // src/ram.vhd(68[19:45])
    defparam i2340_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2339_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_212_3), .O(n2587));   // src/ram.vhd(68[19:45])
    defparam i2339_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2338_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_212_2), .O(n2586));   // src/ram.vhd(68[19:45])
    defparam i2338_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2337_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_212_1), .O(n2585));   // src/ram.vhd(68[19:45])
    defparam i2337_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2336_3_lut_4_lut (.I0(n175), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_212_0), .O(n2584));   // src/ram.vhd(68[19:45])
    defparam i2336_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i176_2_lut_3_lut (.I0(n47), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n176_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i176_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i175_2_lut_3_lut (.I0(n47), .I1(port_id[5]), 
            .I2(port_id[6]), .I3(wea[0]), .O(n175));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i175_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1343_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_87_7), .O(n1591));   // src/ram.vhd(68[19:45])
    defparam i1343_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1342_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_87_6), .O(n1590));   // src/ram.vhd(68[19:45])
    defparam i1342_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1341_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_87_5), .O(n1589));   // src/ram.vhd(68[19:45])
    defparam i1341_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1340_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_87_4), .O(n1588));   // src/ram.vhd(68[19:45])
    defparam i1340_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1339_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_87_3), .O(n1587));   // src/ram.vhd(68[19:45])
    defparam i1339_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1338_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_87_2), .O(n1586));   // src/ram.vhd(68[19:45])
    defparam i1338_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1337_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_87_1), .O(n1585));   // src/ram.vhd(68[19:45])
    defparam i1337_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1336_3_lut_4_lut (.I0(n181), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_87_0), .O(n1584));   // src/ram.vhd(68[19:45])
    defparam i1336_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1335_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[7] ), 
            .I3(ram_s_86_7), .O(n1583));   // src/ram.vhd(68[19:45])
    defparam i1335_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1334_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[6] ), 
            .I3(ram_s_86_6), .O(n1582));   // src/ram.vhd(68[19:45])
    defparam i1334_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i101_2_lut_3_lut_4_lut (.I0(n21), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n101));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i101_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i1333_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[5] ), 
            .I3(ram_s_86_5), .O(n1581));   // src/ram.vhd(68[19:45])
    defparam i1333_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i27_2_lut_3_lut (.I0(n11), .I1(port_id[2]), 
            .I2(port_id[3]), .I3(wea[0]), .O(n27));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i27_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1332_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\sx[4] ), 
            .I3(ram_s_86_4), .O(n1580));   // src/ram.vhd(68[19:45])
    defparam i1332_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1331_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_86_3), .O(n1579));   // src/ram.vhd(68[19:45])
    defparam i1331_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1330_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[10] ), 
            .I3(ram_s_86_2), .O(n1578));   // src/ram.vhd(68[19:45])
    defparam i1330_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1329_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[9] ), 
            .I3(ram_s_86_1), .O(n1577));   // src/ram.vhd(68[19:45])
    defparam i1329_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1328_3_lut_4_lut (.I0(n179), .I1(port_id[7]), .I2(\register_vector[8] ), 
            .I3(ram_s_86_0), .O(n1576));   // src/ram.vhd(68[19:45])
    defparam i1328_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i43_2_lut_3_lut_4_lut (.I0(n11), .I1(port_id[2]), 
            .I2(port_id[3]), .I3(port_id[4]), .O(n43));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i43_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 EnabledDecoder_2_i121_2_lut_3_lut_4_lut (.I0(n18), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n121_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i121_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i123_2_lut_3_lut_4_lut (.I0(n20), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n123_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i123_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i131_2_lut_3_lut_4_lut (.I0(n19), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n131));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i131_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i133_2_lut_3_lut_4_lut (.I0(n21), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n133));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i133_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i100_2_lut_3_lut_4_lut (.I0(n19), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n100));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i100_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i90_2_lut_3_lut_4_lut (.I0(n18), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n90_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i90_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i8316_3_lut (.I0(ram_s_84_6), .I1(ram_s_85_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9375));
    defparam i8316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8317_3_lut (.I0(ram_s_86_6), .I1(ram_s_87_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9376));
    defparam i8317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8293_3_lut (.I0(ram_s_82_6), .I1(ram_s_83_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9352));
    defparam i8293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8292_3_lut (.I0(ram_s_80_6), .I1(ram_s_81_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9351));
    defparam i8292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9045_3_lut (.I0(n14012), .I1(n13916), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10104));
    defparam i9045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9042_3_lut (.I0(n14354), .I1(n14264), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10101));
    defparam i9042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8247_3_lut (.I0(ram_s_68_6), .I1(ram_s_69_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9306));
    defparam i8247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8248_3_lut (.I0(ram_s_70_6), .I1(ram_s_71_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9307));
    defparam i8248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8233_3_lut (.I0(ram_s_66_6), .I1(ram_s_67_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9292));
    defparam i8233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8232_3_lut (.I0(ram_s_64_6), .I1(ram_s_65_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9291));
    defparam i8232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8580_3_lut (.I0(ram_s_148_6), .I1(ram_s_149_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9639));
    defparam i8580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8581_3_lut (.I0(ram_s_150_6), .I1(ram_s_151_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9640));
    defparam i8581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8563_3_lut (.I0(ram_s_146_6), .I1(ram_s_147_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9622));
    defparam i8563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8562_3_lut (.I0(ram_s_144_6), .I1(ram_s_145_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9621));
    defparam i8562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8382_3_lut (.I0(ram_s_100_6), .I1(ram_s_101_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9441));
    defparam i8382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8383_3_lut (.I0(ram_s_102_6), .I1(ram_s_103_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9442));
    defparam i8383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8365_3_lut (.I0(ram_s_98_6), .I1(ram_s_99_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9424));
    defparam i8365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8364_3_lut (.I0(ram_s_96_6), .I1(ram_s_97_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9423));
    defparam i8364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9009_3_lut (.I0(ram_s_244_4), .I1(ram_s_245_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10068));
    defparam i9009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9010_3_lut (.I0(ram_s_246_4), .I1(ram_s_247_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10069));
    defparam i9010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9001_3_lut (.I0(ram_s_242_4), .I1(ram_s_243_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10060));
    defparam i9001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9000_3_lut (.I0(ram_s_240_4), .I1(ram_s_241_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10059));
    defparam i9000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8175_3_lut (.I0(ram_s_52_6), .I1(ram_s_53_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9234));
    defparam i8175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8176_3_lut (.I0(ram_s_54_6), .I1(ram_s_55_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9235));
    defparam i8176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8158_3_lut (.I0(ram_s_50_6), .I1(ram_s_51_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9217));
    defparam i8158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8157_3_lut (.I0(ram_s_48_6), .I1(ram_s_49_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9216));
    defparam i8157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7754_3_lut (.I0(n11324), .I1(n8812), .I2(port_id[3]), .I3(wea[0]), 
            .O(n8813));
    defparam i7754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7753_3_lut (.I0(n12878), .I1(n12812), .I2(port_id[2]), .I3(wea[0]), 
            .O(n8812));
    defparam i7753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7739_3_lut (.I0(n11192), .I1(n13562), .I2(port_id[3]), .I3(wea[0]), 
            .O(n8798));
    defparam i7739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7796_3_lut (.I0(n11516), .I1(n12428), .I2(port_id[3]), .I3(wea[0]), 
            .O(n8855));
    defparam i7796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1259_3_lut_4_lut (.I0(n161), .I1(port_id[7]), .I2(\register_vector[11] ), 
            .I3(ram_s_77_3), .O(n1507));   // src/ram.vhd(68[19:45])
    defparam i1259_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i18_2_lut_4_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[1]), .I3(port_id[2]), .O(n18));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i18_2_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i19_2_lut_4_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[1]), .I3(port_id[2]), .O(n19));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i19_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i17_2_lut_4_lut (.I0(spm_enable), .I1(port_id[0]), 
            .I2(port_id[1]), .I3(port_id[2]), .O(n17));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i17_2_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i9006_3_lut (.I0(ram_s_244_6), .I1(ram_s_245_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10065));
    defparam i9006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9007_3_lut (.I0(ram_s_246_6), .I1(ram_s_247_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10066));
    defparam i9007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8989_3_lut (.I0(ram_s_242_6), .I1(ram_s_243_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10048));
    defparam i8989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8988_3_lut (.I0(ram_s_240_6), .I1(ram_s_241_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10047));
    defparam i8988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8219_3_lut (.I0(n12542), .I1(n9277), .I2(port_id[3]), .I3(wea[0]), 
            .O(n9278));
    defparam i8219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8218_3_lut (.I0(n12638), .I1(n12308), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9277));
    defparam i8218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7766_3_lut (.I0(n11360), .I1(n8824), .I2(port_id[3]), .I3(wea[0]), 
            .O(n8825));
    defparam i7766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7765_3_lut (.I0(n13196), .I1(n13094), .I2(port_id[2]), .I3(wea[0]), 
            .O(n8824));
    defparam i7765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8505_3_lut (.I0(ram_s_12_4), .I1(ram_s_13_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9564));
    defparam i8505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8506_3_lut (.I0(ram_s_14_4), .I1(ram_s_15_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9565));
    defparam i8506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8488_3_lut (.I0(ram_s_10_4), .I1(ram_s_11_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9547));
    defparam i8488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8487_3_lut (.I0(ram_s_8_4), .I1(ram_s_9_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9546));
    defparam i8487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i92_2_lut_3_lut_4_lut (.I0(n20), .I1(port_id[3]), 
            .I2(port_id[4]), .I3(port_id[5]), .O(n92_c));   // src/ram.vhd(68[19:45])
    defparam EnabledDecoder_2_i92_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i8535_3_lut (.I0(ram_s_28_4), .I1(ram_s_29_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9594));
    defparam i8535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8536_3_lut (.I0(ram_s_30_4), .I1(ram_s_31_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9595));
    defparam i8536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8527_3_lut (.I0(ram_s_26_4), .I1(ram_s_27_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9586));
    defparam i8527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8526_3_lut (.I0(ram_s_24_4), .I1(ram_s_25_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9585));
    defparam i8526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7876_3_lut (.I0(n12680), .I1(n12530), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8935));
    defparam i7876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7858_3_lut (.I0(n13532), .I1(n13406), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8917));
    defparam i7858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9882_3_lut (.I0(n13286), .I1(n12488), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10941));
    defparam i9882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9883_3_lut (.I0(n12176), .I1(n11390), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10942));
    defparam i9883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9846_3_lut (.I0(n11672), .I1(n15062), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10905));
    defparam i9846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9822_3_lut (.I0(n11216), .I1(n15128), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10881));
    defparam i9822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9811_3_lut (.I0(n11636), .I1(n11564), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10870));
    defparam i9811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9810_3_lut (.I0(n12344), .I1(n12182), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10869));
    defparam i9810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8655_3_lut (.I0(ram_s_164_6), .I1(ram_s_165_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9714));
    defparam i8655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8656_3_lut (.I0(ram_s_166_6), .I1(ram_s_167_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9715));
    defparam i8656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8635_3_lut (.I0(ram_s_162_6), .I1(ram_s_163_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9694));
    defparam i8635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8634_3_lut (.I0(ram_s_160_6), .I1(ram_s_161_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9693));
    defparam i8634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9756_3_lut (.I0(n15212), .I1(n14030), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10815));
    defparam i9756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9727_3_lut (.I0(n12290), .I1(n11738), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10786));
    defparam i9727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9726_3_lut (.I0(n13646), .I1(n12830), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10785));
    defparam i9726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9753_3_lut (.I0(n12536), .I1(n11582), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10812));
    defparam i9753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9742_3_lut (.I0(n13010), .I1(n12776), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10801));
    defparam i9742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9741_3_lut (.I0(n13622), .I1(n13322), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10800));
    defparam i9741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9687_3_lut (.I0(n14528), .I1(n14216), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10746));
    defparam i9687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9688_3_lut (.I0(n13976), .I1(n13448), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10747));
    defparam i9688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9663_3_lut (.I0(n13136), .I1(n11714), .I2(port_id[2]), .I3(wea[0]), 
            .O(n10722));
    defparam i9663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8922_3_lut (.I0(ram_s_204_5), .I1(ram_s_205_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9981));
    defparam i8922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8923_3_lut (.I0(ram_s_206_5), .I1(ram_s_207_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9982));
    defparam i8923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8854_3_lut (.I0(ram_s_202_5), .I1(ram_s_203_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9913));
    defparam i8854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8853_3_lut (.I0(ram_s_200_5), .I1(ram_s_201_5), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9912));
    defparam i8853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8928_3_lut (.I0(ram_s_204_4), .I1(ram_s_205_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9987));
    defparam i8928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8929_3_lut (.I0(ram_s_206_4), .I1(ram_s_207_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9988));
    defparam i8929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8914_3_lut (.I0(ram_s_202_4), .I1(ram_s_203_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9973));
    defparam i8914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8913_3_lut (.I0(ram_s_200_4), .I1(ram_s_201_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9972));
    defparam i8913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8834_3_lut (.I0(n13940), .I1(n14690), .I2(port_id[5]), .I3(wea[0]), 
            .O(n9893));
    defparam i8834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8395_3_lut (.I0(ram_s_106_6), .I1(ram_s_107_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9454));
    defparam i8395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8394_3_lut (.I0(ram_s_104_6), .I1(ram_s_105_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9453));
    defparam i8394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8421_3_lut (.I0(ram_s_108_6), .I1(ram_s_109_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9480));
    defparam i8421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8422_3_lut (.I0(ram_s_110_6), .I1(ram_s_111_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9481));
    defparam i8422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8873_3_lut (.I0(n14042), .I1(n9931), .I2(port_id[3]), .I3(wea[0]), 
            .O(n9932));
    defparam i8873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8872_3_lut (.I0(n14456), .I1(n14312), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9931));
    defparam i8872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7883_3_lut (.I0(n11792), .I1(n8941), .I2(port_id[5]), .I3(wea[0]), 
            .O(n8942));
    defparam i7883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7882_3_lut (.I0(n12500), .I1(n12314), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8941));
    defparam i7882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7919_3_lut (.I0(n11804), .I1(n8977), .I2(port_id[5]), .I3(wea[0]), 
            .O(n8978));
    defparam i7919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7918_3_lut (.I0(n11402), .I1(n11444), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8977));
    defparam i7918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8950_3_lut (.I0(ram_s_218_4), .I1(ram_s_219_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10009));
    defparam i8950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8949_3_lut (.I0(ram_s_216_4), .I1(ram_s_217_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10008));
    defparam i8949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8958_3_lut (.I0(ram_s_220_4), .I1(ram_s_221_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10017));
    defparam i8958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8959_3_lut (.I0(ram_s_222_4), .I1(ram_s_223_4), .I2(port_id[0]), 
            .I3(wea[0]), .O(n10018));
    defparam i8959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8807_3_lut (.I0(n13868), .I1(n9865), .I2(port_id[3]), .I3(wea[0]), 
            .O(n9866));
    defparam i8807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8806_3_lut (.I0(n14114), .I1(n14066), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9865));
    defparam i8806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8777_3_lut (.I0(n13814), .I1(n9835), .I2(port_id[3]), .I3(wea[0]), 
            .O(n9836));
    defparam i8777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8776_3_lut (.I0(n14708), .I1(n14612), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9835));
    defparam i8776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7745_3_lut (.I0(n11258), .I1(n12974), .I2(port_id[3]), .I3(wea[0]), 
            .O(n8804));
    defparam i7745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8074_3_lut (.I0(ram_s_130_2), .I1(ram_s_131_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9133));
    defparam i8074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8073_3_lut (.I0(ram_s_128_2), .I1(ram_s_129_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9132));
    defparam i8073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8088_3_lut (.I0(ram_s_132_2), .I1(ram_s_133_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9147));
    defparam i8088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8089_3_lut (.I0(ram_s_134_2), .I1(ram_s_135_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9148));
    defparam i8089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8434_3_lut (.I0(ram_s_114_6), .I1(ram_s_115_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9493));
    defparam i8434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8433_3_lut (.I0(ram_s_112_6), .I1(ram_s_113_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9492));
    defparam i8433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8445_3_lut (.I0(ram_s_116_6), .I1(ram_s_117_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9504));
    defparam i8445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8446_3_lut (.I0(ram_s_118_6), .I1(ram_s_119_6), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9505));
    defparam i8446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8065_3_lut (.I0(ram_s_10_7), .I1(ram_s_11_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9124));
    defparam i8065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8064_3_lut (.I0(ram_s_8_7), .I1(ram_s_9_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9123));
    defparam i8064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8097_3_lut (.I0(ram_s_12_7), .I1(ram_s_13_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9156));
    defparam i8097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8098_3_lut (.I0(ram_s_14_7), .I1(ram_s_15_7), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9157));
    defparam i8098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8143_3_lut (.I0(ram_s_146_2), .I1(ram_s_147_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9202));
    defparam i8143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8142_3_lut (.I0(ram_s_144_2), .I1(ram_s_145_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9201));
    defparam i8142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8154_3_lut (.I0(ram_s_148_2), .I1(ram_s_149_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9213));
    defparam i8154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8155_3_lut (.I0(ram_s_150_2), .I1(ram_s_151_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9214));
    defparam i8155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7789_3_lut (.I0(n12560), .I1(n11702), .I2(port_id[2]), .I3(wea[0]), 
            .O(n8848));
    defparam i7789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8428_3_lut (.I0(ram_s_210_2), .I1(ram_s_211_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9487));
    defparam i8428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8427_3_lut (.I0(ram_s_208_2), .I1(ram_s_209_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9486));
    defparam i8427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8439_3_lut (.I0(ram_s_212_2), .I1(ram_s_213_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9498));
    defparam i8439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8440_3_lut (.I0(ram_s_214_2), .I1(ram_s_215_2), .I2(port_id[0]), 
            .I3(wea[0]), .O(n9499));
    defparam i8440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7894_3_lut (.I0(n12230), .I1(n12080), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8953));
    defparam i7894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7911_3_lut (.I0(n12020), .I1(n11570), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8970));
    defparam i7911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7912_3_lut (.I0(n11420), .I1(n11972), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8971));
    defparam i7912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7982_3_lut (.I0(n11852), .I1(n9040), .I2(port_id[3]), .I3(wea[0]), 
            .O(n9041));
    defparam i7982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7981_3_lut (.I0(n12848), .I1(n11870), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9040));
    defparam i7981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8442_3_lut (.I0(n11684), .I1(n11246), .I2(port_id[4]), .I3(wea[0]), 
            .O(n9501));
    defparam i8442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8413_3_lut (.I0(n13592), .I1(n13478), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9472));
    defparam i8413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8416_3_lut (.I0(n13328), .I1(n13190), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9475));
    defparam i8416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8788_3_lut (.I0(n14414), .I1(n14276), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9847));
    defparam i8788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8371_3_lut (.I0(n14930), .I1(n14804), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9430));
    defparam i8371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8374_3_lut (.I0(n14684), .I1(n14552), .I2(port_id[2]), .I3(wea[0]), 
            .O(n9433));
    defparam i8374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7784_3_lut (.I0(n11462), .I1(n8842), .I2(port_id[5]), .I3(wea[0]), 
            .O(n8843));
    defparam i7784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7783_3_lut (.I0(n12590), .I1(n11888), .I2(port_id[4]), .I3(wea[0]), 
            .O(n8842));
    defparam i7783_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module shift_and_rotate_operations
//

module shift_and_rotate_operations (shift_rotate_result, CLK_3P3_MHZ_c, 
            \instruction[7] , \sx[6] , \instruction[3] , wea, \sx[5] , 
            \sx[7] , \sx[4] , \register_vector[11] , \register_vector[10] , 
            \register_vector[9] , \register_vector[8] , \instruction[2] , 
            \instruction[0] , \instruction[1] , carry_flag);
    output [7:0]shift_rotate_result;
    input CLK_3P3_MHZ_c;
    input \instruction[7] ;
    input \sx[6] ;
    input \instruction[3] ;
    input [0:0]wea;
    input \sx[5] ;
    input \sx[7] ;
    input \sx[4] ;
    input \register_vector[11] ;
    input \register_vector[10] ;
    input \register_vector[9] ;
    input \register_vector[8] ;
    input \instruction[2] ;
    input \instruction[0] ;
    input \instruction[1] ;
    input carry_flag;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [7:0]shift_rotate_value;   // src/shift_and_rotate_operations.vhd(47[12:30])
    
    wire shift_in_bit, n12503;
    
    SB_DFFSS shift_rotate_result_i0 (.Q(shift_rotate_result[0]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[0]), .S(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_DFFSR shift_rotate_result_i1 (.Q(shift_rotate_result[1]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[1]), .R(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_DFFSR shift_rotate_result_i2 (.Q(shift_rotate_result[2]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[2]), .R(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_DFFSR shift_rotate_result_i3 (.Q(shift_rotate_result[3]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[3]), .R(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_DFFSR shift_rotate_result_i4 (.Q(shift_rotate_result[4]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[4]), .R(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_DFFSR shift_rotate_result_i5 (.Q(shift_rotate_result[5]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[5]), .R(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_DFFSS shift_rotate_result_i6 (.Q(shift_rotate_result[6]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[6]), .S(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_DFFSR shift_rotate_result_i7 (.Q(shift_rotate_result[7]), .C(CLK_3P3_MHZ_c), 
            .D(shift_rotate_value[7]), .R(\instruction[7] ));   // src/shift_and_rotate_operations.vhd(53[9] 59[16])
    SB_LUT4 i36_3_lut (.I0(\sx[6] ), .I1(shift_in_bit), .I2(\instruction[3] ), 
            .I3(wea[0]), .O(shift_rotate_value[7]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35_3_lut (.I0(\sx[5] ), .I1(\sx[7] ), .I2(\instruction[3] ), 
            .I3(wea[0]), .O(shift_rotate_value[6]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i35_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34_3_lut (.I0(\sx[4] ), .I1(\sx[6] ), .I2(\instruction[3] ), 
            .I3(wea[0]), .O(shift_rotate_value[5]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut (.I0(\register_vector[11] ), .I1(\sx[5] ), .I2(\instruction[3] ), 
            .I3(wea[0]), .O(shift_rotate_value[4]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i33_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32_3_lut (.I0(\register_vector[10] ), .I1(\sx[4] ), .I2(\instruction[3] ), 
            .I3(wea[0]), .O(shift_rotate_value[3]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31_3_lut (.I0(\register_vector[9] ), .I1(\register_vector[11] ), 
            .I2(\instruction[3] ), .I3(wea[0]), .O(shift_rotate_value[2]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30_3_lut (.I0(\register_vector[8] ), .I1(\register_vector[10] ), 
            .I2(\instruction[3] ), .I3(wea[0]), .O(shift_rotate_value[1]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut (.I0(shift_in_bit), .I1(\register_vector[9] ), .I2(\instruction[3] ), 
            .I3(wea[0]), .O(shift_rotate_value[0]));   // src/shift_and_rotate_operations.vhd(170[13] 171[57])
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 instruction_2__bdd_4_lut (.I0(\instruction[2] ), .I1(\sx[7] ), 
            .I2(\instruction[0] ), .I3(\instruction[1] ), .O(n12503));
    defparam instruction_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12503_bdd_4_lut (.I0(n12503), .I1(\register_vector[8] ), .I2(carry_flag), 
            .I3(\instruction[1] ), .O(shift_in_bit));
    defparam n12503_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module sel_of_out_port_value
//

module sel_of_out_port_value (\register_vector[8] , \instruction[4] , \instruction[13] , 
            LED1_c_0, wea);
    input \register_vector[8] ;
    input \instruction[4] ;
    input \instruction[13] ;
    output LED1_c_0;
    input [0:0]wea;
    
    
    SB_LUT4 i10_3_lut (.I0(\register_vector[8] ), .I1(\instruction[4] ), 
            .I2(\instruction[13] ), .I3(wea[0]), .O(LED1_c_0));   // src/sel_of_out_port_value.vhd(140[14] 141[62])
    defparam i10_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module sel_of_2nd_op_to_alu_and_port_id
//

module sel_of_2nd_op_to_alu_and_port_id (\register_vector[7] , \instruction[7] , 
            \instruction[12] , port_id, wea, \register_vector[2] , \instruction[2] , 
            \register_vector[3] , \instruction[3] , \register_vector[4] , 
            \instruction[4] , \register_vector[6] , \instruction[6] , 
            \register_vector[5] , \instruction[5] , \register_vector[1] , 
            \instruction[1] , \register_vector[0] , \instruction[0] );
    input \register_vector[7] ;
    input \instruction[7] ;
    input \instruction[12] ;
    output [7:0]port_id;
    input [0:0]wea;
    input \register_vector[2] ;
    input \instruction[2] ;
    input \register_vector[3] ;
    input \instruction[3] ;
    input \register_vector[4] ;
    input \instruction[4] ;
    input \register_vector[6] ;
    input \instruction[6] ;
    input \register_vector[5] ;
    input \instruction[5] ;
    input \register_vector[1] ;
    input \instruction[1] ;
    input \register_vector[0] ;
    input \instruction[0] ;
    
    
    SB_LUT4 i29_3_lut (.I0(\register_vector[7] ), .I1(\instruction[7] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[7]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut (.I0(\register_vector[2] ), .I1(\instruction[2] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[2]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_3_lut (.I0(\register_vector[3] ), .I1(\instruction[3] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[3]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26_3_lut (.I0(\register_vector[4] ), .I1(\instruction[4] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[4]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28_3_lut (.I0(\register_vector[6] ), .I1(\instruction[6] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[6]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27_3_lut (.I0(\register_vector[5] ), .I1(\instruction[5] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[5]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_3_lut (.I0(\register_vector[1] ), .I1(\instruction[1] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[1]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_3_lut (.I0(\register_vector[0] ), .I1(\instruction[0] ), 
            .I2(\instruction[12] ), .I3(wea[0]), .O(port_id[0]));   // src/sel_of_2nd_op_to_alu_and_port_id.vhd(141[14] 142[60])
    defparam i9_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module register_bank_control
//

module register_bank_control (sx_addr4_value, \sx_addr[4] , CLK_3P3_MHZ_c, 
            internal_reset_N_50, \sy_addr[4] , flag_enable_type_N_217, 
            \instruction[16] , \instruction[14] , \instruction[17] , loadstar_type, 
            regbank_type_N_77, \instruction[15] , n4283, wea, \instruction[12] , 
            \t_state[1] , shadow_bank, \instruction[0] , internal_reset);
    input sx_addr4_value;
    output \sx_addr[4] ;
    input CLK_3P3_MHZ_c;
    input internal_reset_N_50;
    output \sy_addr[4] ;
    input flag_enable_type_N_217;
    input \instruction[16] ;
    input \instruction[14] ;
    input \instruction[17] ;
    output loadstar_type;
    output regbank_type_N_77;
    input \instruction[15] ;
    input n4283;
    input [0:0]wea;
    input \instruction[12] ;
    input \t_state[1] ;
    input shadow_bank;
    input \instruction[0] ;
    input internal_reset;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    wire bank_value_N_92, n8744, regbank_type_N_85, regbank_type_N_74, 
        n6, n758;
    
    SB_DFF sx_addr_4_43 (.Q(\sx_addr[4] ), .C(CLK_3P3_MHZ_c), .D(sx_addr4_value));   // src/register_bank_control.vhd(57[9] 59[16])
    SB_DFFESS bank_44 (.Q(\sy_addr[4] ), .C(CLK_3P3_MHZ_c), .E(internal_reset_N_50), 
            .D(bank_value_N_92), .S(n8744));   // src/register_bank_control.vhd(63[9] 67[16])
    SB_LUT4 i1_2_lut_4_lut (.I0(flag_enable_type_N_217), .I1(\instruction[16] ), 
            .I2(\instruction[14] ), .I3(\instruction[17] ), .O(regbank_type_N_85));   // src/register_bank_control.vhd(81[7] 82[69])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut_adj_297 (.I0(flag_enable_type_N_217), .I1(\instruction[16] ), 
            .I2(\instruction[14] ), .I3(\instruction[17] ), .O(loadstar_type));   // src/register_bank_control.vhd(81[7] 82[69])
    defparam i1_2_lut_4_lut_adj_297.LUT_INIT = 16'h0080;
    SB_LUT4 i2_3_lut (.I0(regbank_type_N_77), .I1(\instruction[15] ), .I2(n4283), 
            .I3(wea[0]), .O(regbank_type_N_74));   // src/register_bank_control.vhd(79[19] 80[77])
    defparam i2_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i2_4_lut (.I0(\instruction[12] ), .I1(\t_state[1] ), .I2(regbank_type_N_74), 
            .I3(regbank_type_N_85), .O(n6));   // src/register_bank_control.vhd(63[9] 67[16])
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i611_3_lut (.I0(shadow_bank), .I1(\instruction[0] ), .I2(\instruction[16] ), 
            .I3(wea[0]), .O(n758));   // src/register_bank_control.vhd(93[16] 96[85])
    defparam i611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i79_2_lut (.I0(\sy_addr[4] ), .I1(n6), .I2(wea[0]), .I3(wea[0]), 
            .O(bank_value_N_92));   // src/register_bank_control.vhd(93[16] 94[34])
    defparam i79_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 instruction_17_downto_4_17__I_0_45_2_lut (.I0(\instruction[17] ), 
            .I1(\instruction[16] ), .I2(wea[0]), .I3(wea[0]), .O(regbank_type_N_77));   // src/register_bank_control.vhd(79[19:82])
    defparam instruction_17_downto_4_17__I_0_45_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_3_lut_3_lut (.I0(internal_reset), .I1(n6), .I2(n758), .I3(wea[0]), 
            .O(n8744));   // src/register_bank_control.vhd(63[9] 67[16])
    defparam i3_3_lut_3_lut.LUT_INIT = 16'h4040;
    
endmodule
//
// Verilog Description of module program_counter
//

module program_counter (n765, address, CLK_3P3_MHZ_c, internal_reset, 
            n938, \pc_mode[0] , wea, \pc_value[0] , \pc_vector[1] , 
            register_vector, \instruction[0] , \return_vector[0] , \instruction[12] , 
            \pc_vector[2] , \pc_mode_2__N_158[2] , pc_mode_2__N_104, \instruction[3] , 
            \return_vector[3] , \instruction[17] , \instruction[16] , 
            n6, \pc_vector[4] , \pc_vector[5] , \pc_vector[6] , \pc_vector[11] , 
            \pc_vector[10] , \instruction[9] , \return_vector[9] , \pc_vector[8] , 
            \pc_vector[7] );
    input n765;
    output [11:0]address;
    input CLK_3P3_MHZ_c;
    input internal_reset;
    input n938;
    input \pc_mode[0] ;
    input [0:0]wea;
    output \pc_value[0] ;
    input \pc_vector[1] ;
    input [11:0]register_vector;
    input \instruction[0] ;
    input \return_vector[0] ;
    input \instruction[12] ;
    input \pc_vector[2] ;
    input \pc_mode_2__N_158[2] ;
    input pc_mode_2__N_104;
    input \instruction[3] ;
    input \return_vector[3] ;
    input \instruction[17] ;
    input \instruction[16] ;
    input n6;
    input \pc_vector[4] ;
    input \pc_vector[5] ;
    input \pc_vector[6] ;
    input \pc_vector[11] ;
    input \pc_vector[10] ;
    input \instruction[9] ;
    input \return_vector[9] ;
    input \pc_vector[8] ;
    input \pc_vector[7] ;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [11:0]pc_value;   // src/program_counter.vhd(48[12:20])
    
    wire n232;
    wire [11:0]half_pc;   // src/program_counter.vhd(49[12:19])
    
    wire n223, n229, n217, pc_value_0__N_530, pc_value_0__N_520, n6_c, 
        pc_value_0__N_513;
    wire [10:0]half_pc_11__N_591;
    
    wire n5, n6_adj_817, n6_adj_818;
    wire [10:0]n317;
    
    wire n6_adj_819, n6_adj_821, n6_adj_822, n6_adj_823, n6_adj_824, 
        n238, n6_adj_825, n6_adj_826, n6_adj_828, n6_adj_829;
    
    SB_DFFESR pc__i5 (.Q(address[5]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[5]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i4 (.Q(address[4]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[4]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i3 (.Q(address[3]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[3]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i2 (.Q(address[2]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[2]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i1 (.Q(address[1]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[1]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFF pc__i0 (.Q(address[0]), .C(CLK_3P3_MHZ_c), .D(n938));   // src/program_counter.vhd(55[9] 61[16])
    SB_LUT4 half_pc_11__I_0_i9_3_lut_4_lut (.I0(n232), .I1(half_pc[8]), 
            .I2(\pc_mode[0] ), .I3(half_pc[9]), .O(pc_value[9]));   // src/program_counter.vhd(367[9] 374[18])
    defparam half_pc_11__I_0_i9_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i106_2_lut_3_lut (.I0(n223), .I1(half_pc[5]), .I2(half_pc[6]), 
            .I3(wea[0]), .O(n229));   // src/program_counter.vhd(328[9] 335[18])
    defparam i106_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 half_pc_11__I_0_i6_3_lut_4_lut (.I0(n223), .I1(half_pc[5]), 
            .I2(\pc_mode[0] ), .I3(half_pc[6]), .O(pc_value[6]));   // src/program_counter.vhd(328[9] 335[18])
    defparam half_pc_11__I_0_i6_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_DFFESR pc__i6 (.Q(address[6]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[6]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_LUT4 half_pc_11__I_0_i4_3_lut_4_lut (.I0(n217), .I1(half_pc[3]), 
            .I2(\pc_mode[0] ), .I3(half_pc[4]), .O(pc_value[4]));   // src/program_counter.vhd(302[9] 309[18])
    defparam half_pc_11__I_0_i4_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i100_2_lut_3_lut (.I0(n217), .I1(half_pc[3]), .I2(half_pc[4]), 
            .I3(wea[0]), .O(n223));   // src/program_counter.vhd(302[9] 309[18])
    defparam i100_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 half_pc_11__I_0_i2_3_lut_4_lut (.I0(\pc_value[0] ), .I1(half_pc[1]), 
            .I2(\pc_mode[0] ), .I3(half_pc[2]), .O(pc_value[2]));   // src/program_counter.vhd(276[9] 283[18])
    defparam half_pc_11__I_0_i2_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i94_2_lut_3_lut (.I0(\pc_value[0] ), .I1(half_pc[1]), .I2(half_pc[2]), 
            .I3(wea[0]), .O(n217));   // src/program_counter.vhd(276[9] 283[18])
    defparam i94_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 half_pc_11__I_0_i1_3_lut (.I0(half_pc[1]), .I1(\pc_mode[0] ), 
            .I2(\pc_value[0] ), .I3(wea[0]), .O(pc_value[1]));   // src/program_counter.vhd(258[21:49])
    defparam half_pc_11__I_0_i1_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 half_pc_11__I_0_i3_3_lut (.I0(half_pc[3]), .I1(\pc_mode[0] ), 
            .I2(n217), .I3(wea[0]), .O(pc_value[3]));   // src/program_counter.vhd(258[21:49])
    defparam half_pc_11__I_0_i3_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 i2_4_lut (.I0(pc_value_0__N_530), .I1(pc_value_0__N_520), .I2(\pc_vector[1] ), 
            .I3(register_vector[1]), .O(n6_c));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut (.I0(pc_value_0__N_513), .I1(n6_c), .I2(half_pc_11__N_591[10]), 
            .I3(address[1]), .O(half_pc[1]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i612_4_lut (.I0(\instruction[0] ), .I1(\pc_mode[0] ), .I2(\return_vector[0] ), 
            .I3(\instruction[12] ), .O(n5));   // src/program_counter.vhd(76[4] 80[71])
    defparam i612_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i2_4_lut_adj_276 (.I0(pc_value_0__N_530), .I1(half_pc_11__N_591[10]), 
            .I2(n5), .I3(address[0]), .O(n6_adj_817));   // src/program_counter.vhd(76[4] 80[71])
    defparam i2_4_lut_adj_276.LUT_INIT = 16'ha0ec;
    SB_LUT4 i3_4_lut_adj_277 (.I0(pc_value_0__N_513), .I1(n6_adj_817), .I2(pc_value_0__N_520), 
            .I3(register_vector[0]), .O(\pc_value[0] ));   // src/program_counter.vhd(76[4] 80[71])
    defparam i3_4_lut_adj_277.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_4_lut_adj_278 (.I0(half_pc_11__N_591[10]), .I1(pc_value_0__N_520), 
            .I2(address[2]), .I3(register_vector[2]), .O(n6_adj_818));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_278.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_279 (.I0(pc_value_0__N_513), .I1(n6_adj_818), .I2(pc_value_0__N_530), 
            .I3(\pc_vector[2] ), .O(half_pc[2]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_279.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_3_lut (.I0(\pc_mode_2__N_158[2] ), .I1(\pc_mode[0] ), .I2(pc_mode_2__N_104), 
            .I3(wea[0]), .O(half_pc_11__N_591[10]));
    defparam i2_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 and_274_i11_2_lut (.I0(\pc_mode_2__N_158[2] ), .I1(\pc_mode[0] ), 
            .I2(wea[0]), .I3(wea[0]), .O(pc_value_0__N_520));   // src/program_counter.vhd(244[5:34])
    defparam and_274_i11_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 and_270_i3_4_lut (.I0(pc_value_0__N_530), .I1(\instruction[3] ), 
            .I2(\return_vector[3] ), .I3(\instruction[12] ), .O(n317[2]));   // src/program_counter.vhd(242[5:52])
    defparam and_270_i3_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i3_4_lut_adj_280 (.I0(n317[2]), .I1(n6_adj_819), .I2(half_pc_11__N_591[10]), 
            .I3(address[3]), .O(half_pc[3]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_280.LUT_INIT = 16'hfeee;
    SB_LUT4 and_269_i11_2_lut (.I0(\pc_mode_2__N_158[2] ), .I1(pc_mode_2__N_104), 
            .I2(wea[0]), .I3(wea[0]), .O(pc_value_0__N_530));   // src/program_counter.vhd(242[5:34])
    defparam and_269_i11_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4_4_lut (.I0(\instruction[17] ), .I1(\pc_mode[0] ), .I2(\instruction[16] ), 
            .I3(n6), .O(pc_value_0__N_513));   // src/program_counter.vhd(243[5:53])
    defparam i4_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i2_4_lut_adj_281 (.I0(half_pc_11__N_591[10]), .I1(pc_value_0__N_520), 
            .I2(address[4]), .I3(register_vector[4]), .O(n6_adj_821));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_281.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_282 (.I0(pc_value_0__N_513), .I1(n6_adj_821), .I2(pc_value_0__N_530), 
            .I3(\pc_vector[4] ), .O(half_pc[4]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_282.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_4_lut_adj_283 (.I0(pc_value_0__N_530), .I1(pc_value_0__N_520), 
            .I2(\pc_vector[5] ), .I3(register_vector[5]), .O(n6_adj_822));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_283.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_284 (.I0(pc_value_0__N_513), .I1(n6_adj_822), .I2(half_pc_11__N_591[10]), 
            .I3(address[5]), .O(half_pc[5]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_284.LUT_INIT = 16'hfeee;
    SB_LUT4 half_pc_11__I_0_i5_3_lut (.I0(half_pc[5]), .I1(\pc_mode[0] ), 
            .I2(n223), .I3(wea[0]), .O(pc_value[5]));   // src/program_counter.vhd(258[21:49])
    defparam half_pc_11__I_0_i5_3_lut.LUT_INIT = 16'ha6a6;
    SB_DFFESR pc__i11 (.Q(address[11]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[11]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i10 (.Q(address[10]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[10]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i9 (.Q(address[9]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[9]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i8 (.Q(address[8]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[8]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_DFFESR pc__i7 (.Q(address[7]), .C(CLK_3P3_MHZ_c), .E(n765), .D(pc_value[7]), 
            .R(internal_reset));   // src/program_counter.vhd(55[9] 61[16])
    SB_LUT4 half_pc_11__I_0_i8_3_lut_4_lut (.I0(half_pc[8]), .I1(\pc_mode[0] ), 
            .I2(n229), .I3(half_pc[7]), .O(pc_value[8]));   // src/program_counter.vhd(258[21:49])
    defparam half_pc_11__I_0_i8_3_lut_4_lut.LUT_INIT = 16'ha6aa;
    SB_LUT4 i2_3_lut_4_lut (.I0(pc_value_0__N_513), .I1(\pc_mode_2__N_158[2] ), 
            .I2(\pc_mode[0] ), .I3(register_vector[9]), .O(n6_adj_823));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'haeaa;
    SB_LUT4 i2_3_lut_4_lut_adj_285 (.I0(pc_value_0__N_513), .I1(\pc_mode_2__N_158[2] ), 
            .I2(\pc_mode[0] ), .I3(register_vector[3]), .O(n6_adj_819));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_3_lut_4_lut_adj_285.LUT_INIT = 16'haeaa;
    SB_LUT4 i3_4_lut_adj_286 (.I0(pc_value_0__N_513), .I1(n6_adj_824), .I2(half_pc_11__N_591[10]), 
            .I3(address[6]), .O(half_pc[6]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_286.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_4_lut_adj_287 (.I0(pc_value_0__N_520), .I1(pc_value_0__N_530), 
            .I2(register_vector[6]), .I3(\pc_vector[6] ), .O(n6_adj_824));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_287.LUT_INIT = 16'heca0;
    SB_LUT4 half_pc_11__I_0_i11_4_lut (.I0(half_pc[11]), .I1(n238), .I2(half_pc[10]), 
            .I3(\pc_mode[0] ), .O(pc_value[11]));   // src/program_counter.vhd(258[21:49])
    defparam half_pc_11__I_0_i11_4_lut.LUT_INIT = 16'h9aaa;
    SB_LUT4 i3_4_lut_adj_288 (.I0(pc_value_0__N_513), .I1(n6_adj_825), .I2(half_pc_11__N_591[10]), 
            .I3(address[11]), .O(half_pc[11]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_288.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_4_lut_adj_289 (.I0(pc_value_0__N_530), .I1(pc_value_0__N_520), 
            .I2(\pc_vector[11] ), .I3(register_vector[11]), .O(n6_adj_825));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_289.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_290 (.I0(pc_value_0__N_513), .I1(n6_adj_826), .I2(half_pc_11__N_591[10]), 
            .I3(address[10]), .O(half_pc[10]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_290.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_4_lut_adj_291 (.I0(pc_value_0__N_520), .I1(pc_value_0__N_530), 
            .I2(register_vector[10]), .I3(\pc_vector[10] ), .O(n6_adj_826));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_291.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_292 (.I0(n317[8]), .I1(n6_adj_823), .I2(half_pc_11__N_591[10]), 
            .I3(address[9]), .O(half_pc[9]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_292.LUT_INIT = 16'hfeee;
    SB_LUT4 and_270_i9_4_lut (.I0(pc_value_0__N_530), .I1(\instruction[9] ), 
            .I2(\return_vector[9] ), .I3(\instruction[12] ), .O(n317[8]));   // src/program_counter.vhd(242[5:52])
    defparam and_270_i9_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i109_2_lut (.I0(n229), .I1(half_pc[7]), .I2(wea[0]), .I3(wea[0]), 
            .O(n232));   // src/program_counter.vhd(354[9] 361[18])
    defparam i109_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_293 (.I0(pc_value_0__N_513), .I1(n6_adj_828), .I2(half_pc_11__N_591[10]), 
            .I3(address[8]), .O(half_pc[8]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_293.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_4_lut_adj_294 (.I0(pc_value_0__N_520), .I1(pc_value_0__N_530), 
            .I2(register_vector[8]), .I3(\pc_vector[8] ), .O(n6_adj_828));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_294.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_295 (.I0(pc_value_0__N_513), .I1(n6_adj_829), .I2(half_pc_11__N_591[10]), 
            .I3(address[7]), .O(half_pc[7]));   // src/program_counter.vhd(242[4] 245[65])
    defparam i3_4_lut_adj_295.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_4_lut_adj_296 (.I0(pc_value_0__N_530), .I1(pc_value_0__N_520), 
            .I2(\pc_vector[7] ), .I3(register_vector[7]), .O(n6_adj_829));   // src/program_counter.vhd(242[4] 245[65])
    defparam i2_4_lut_adj_296.LUT_INIT = 16'heca0;
    SB_LUT4 half_pc_11__I_0_i10_3_lut (.I0(half_pc[10]), .I1(\pc_mode[0] ), 
            .I2(n238), .I3(wea[0]), .O(pc_value[10]));   // src/program_counter.vhd(258[21:49])
    defparam half_pc_11__I_0_i10_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 half_pc_11__I_0_i7_3_lut (.I0(half_pc[7]), .I1(\pc_mode[0] ), 
            .I2(n229), .I3(wea[0]), .O(pc_value[7]));   // src/program_counter.vhd(258[21:49])
    defparam half_pc_11__I_0_i7_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 i115_2_lut_3_lut_4_lut (.I0(n229), .I1(half_pc[7]), .I2(half_pc[8]), 
            .I3(half_pc[9]), .O(n238));   // src/program_counter.vhd(367[9] 374[18])
    defparam i115_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    
endmodule
//
// Verilog Description of module mux_outputs_from_alu_spm_input_ports
//

module mux_outputs_from_alu_spm_input_ports (arith_logical_result, shift_rotate_result, 
            alu_mux_sel, wea, spm_data, alu_result);
    input [7:0]arith_logical_result;
    input [7:0]shift_rotate_result;
    input [1:0]alu_mux_sel;
    input [0:0]wea;
    input [7:0]spm_data;
    output [7:0]alu_result;
    
    
    wire n1, n1_adj_810, n1_adj_811, n1_adj_812, n1_adj_813, n1_adj_814, 
        n1_adj_815, n1_adj_816;
    
    SB_LUT4 alu_mux_sel_1__I_0_Mux_0_i1_3_lut (.I0(arith_logical_result[0]), 
            .I1(shift_rotate_result[0]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_0_i3_4_lut (.I0(n1), .I1(spm_data[0]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[0]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_0_i3_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_1_i1_3_lut (.I0(arith_logical_result[1]), 
            .I1(shift_rotate_result[1]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1_adj_810));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_1_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_1_i3_4_lut (.I0(n1_adj_810), .I1(spm_data[1]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[1]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_1_i3_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_2_i1_3_lut (.I0(arith_logical_result[2]), 
            .I1(shift_rotate_result[2]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1_adj_811));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_2_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_2_i3_4_lut (.I0(n1_adj_811), .I1(spm_data[2]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[2]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_2_i3_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_3_i1_3_lut (.I0(arith_logical_result[3]), 
            .I1(shift_rotate_result[3]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1_adj_812));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_3_i3_4_lut (.I0(n1_adj_812), .I1(spm_data[3]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[3]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_3_i3_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_4_i1_3_lut (.I0(arith_logical_result[4]), 
            .I1(shift_rotate_result[4]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1_adj_813));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_4_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_4_i3_4_lut (.I0(n1_adj_813), .I1(spm_data[4]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[4]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_4_i3_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_5_i1_3_lut (.I0(arith_logical_result[5]), 
            .I1(shift_rotate_result[5]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1_adj_814));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_5_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_5_i3_4_lut (.I0(n1_adj_814), .I1(spm_data[5]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[5]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_5_i3_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_6_i1_3_lut (.I0(arith_logical_result[6]), 
            .I1(shift_rotate_result[6]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1_adj_815));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_6_i3_4_lut (.I0(n1_adj_815), .I1(spm_data[6]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[6]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_6_i3_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_7_i1_3_lut (.I0(arith_logical_result[7]), 
            .I1(shift_rotate_result[7]), .I2(alu_mux_sel[0]), .I3(wea[0]), 
            .O(n1_adj_816));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_7_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 alu_mux_sel_1__I_0_Mux_7_i3_4_lut (.I0(n1_adj_816), .I1(spm_data[7]), 
            .I2(alu_mux_sel[1]), .I3(alu_mux_sel[0]), .O(alu_result[7]));   // src/mux_outputs_from_alu_spm_input_ports.vhd(52[9] 63[18])
    defparam alu_mux_sel_1__I_0_Mux_7_i3_4_lut.LUT_INIT = 16'hca0a;
    
endmodule
//
// Verilog Description of module flags
//

module flags (CLK_3P3_MHZ_c, instruction_13_N_701, carry_arith_logical_7, 
            zero_flag, internal_reset, carry_flag, \instruction[13] , 
            carry_flag_value_N_436, flag_enable_type_N_216, arith_carry_in, 
            arith_logical_result, wea, \alu_mux_sel_value[1] , alu_mux_sel_value_0__N_184, 
            \instruction[14] , arith_logical_sel_2__N_179, flag_enable, 
            alu_result, \instruction[15] , \instruction[16] , shadow_zero_flag, 
            \arith_logical_sel[0] , \arith_logical_sel[2] , n11080, \register_vector[9] , 
            n338, n3783, n4, n11084, \port_id[1] , \half_arith_logical[1] , 
            \sx[7] , \register_vector[8] , \instruction[3] , shadow_carry_flag, 
            \instruction[7] , \port_id[5] , n722, n11107, \sx[5] , 
            n11109, n350, \half_arith_logical[5] , n4_adj_2);
    input CLK_3P3_MHZ_c;
    input instruction_13_N_701;
    input carry_arith_logical_7;
    output zero_flag;
    input internal_reset;
    output carry_flag;
    input \instruction[13] ;
    input carry_flag_value_N_436;
    input flag_enable_type_N_216;
    output arith_carry_in;
    input [7:0]arith_logical_result;
    input [0:0]wea;
    input \alu_mux_sel_value[1] ;
    input alu_mux_sel_value_0__N_184;
    input \instruction[14] ;
    input arith_logical_sel_2__N_179;
    input flag_enable;
    input [7:0]alu_result;
    input \instruction[15] ;
    input \instruction[16] ;
    input shadow_zero_flag;
    output \arith_logical_sel[0] ;
    input \arith_logical_sel[2] ;
    input n11080;
    input \register_vector[9] ;
    input n338;
    output n3783;
    input n4;
    output n11084;
    input \port_id[1] ;
    output \half_arith_logical[1] ;
    input \sx[7] ;
    input \register_vector[8] ;
    input \instruction[3] ;
    input shadow_carry_flag;
    input \instruction[7] ;
    input \port_id[5] ;
    input n722;
    input n11107;
    input \sx[5] ;
    input n11109;
    input n350;
    output \half_arith_logical[5] ;
    output n4_adj_2;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    wire shift_carry_value_N_413, shift_carry, n687, n207, use_zero_flag, 
        arith_carry, zero_flag_value, n761, carry_flag_value, lower_parity, 
        n55, n8728, n4_c, n4_adj_806, n8718, parity, n5, n4_adj_807, 
        n8787, n8783, n8791, upper_zero_sel, n11087, n11163, n7, 
        n12779;
    
    SB_DFFSS shift_carry_423 (.Q(shift_carry), .C(CLK_3P3_MHZ_c), .D(shift_carry_value_N_413), 
            .S(n687));   // src/flags.vhd(83[9] 87[16])
    SB_DFFSR use_zero_flag_424 (.Q(use_zero_flag), .C(CLK_3P3_MHZ_c), .D(n207), 
            .R(instruction_13_N_701));   // src/flags.vhd(83[9] 87[16])
    SB_DFF arith_carry_422 (.Q(arith_carry), .C(CLK_3P3_MHZ_c), .D(carry_arith_logical_7));   // src/flags.vhd(83[9] 87[16])
    SB_DFFESR zero_flag_425 (.Q(zero_flag), .C(CLK_3P3_MHZ_c), .E(n761), 
            .D(zero_flag_value), .R(internal_reset));   // src/flags.vhd(91[9] 99[16])
    SB_DFFESR carry_flag_426 (.Q(carry_flag), .C(CLK_3P3_MHZ_c), .E(n761), 
            .D(carry_flag_value), .R(internal_reset));   // src/flags.vhd(91[9] 99[16])
    SB_LUT4 i10092_3_lut_4_lut (.I0(carry_flag), .I1(\instruction[13] ), 
            .I2(carry_flag_value_N_436), .I3(flag_enable_type_N_216), .O(arith_carry_in));
    defparam i10092_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i30_3_lut_4_lut (.I0(carry_flag), .I1(\instruction[13] ), .I2(arith_logical_result[1]), 
            .I3(arith_logical_result[0]), .O(lower_parity));
    defparam i30_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i159_2_lut (.I0(arith_logical_result[3]), .I1(arith_logical_result[2]), 
            .I2(wea[0]), .I3(wea[0]), .O(n55));   // src/flags.vhd(147[9] 148[194])
    defparam i159_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n55), .I1(arith_logical_result[5]), .I2(n8728), 
            .I3(n4_c), .O(n4_adj_806));   // src/flags.vhd(147[9] 178[178])
    defparam i1_4_lut.LUT_INIT = 16'h7350;
    SB_LUT4 lower_parity_I_0_4_lut (.I0(lower_parity), .I1(n55), .I2(n4_adj_806), 
            .I3(n8718), .O(parity));   // src/flags.vhd(106[15:50])
    defparam lower_parity_I_0_4_lut.LUT_INIT = 16'h565a;
    SB_LUT4 i1_4_lut_adj_273 (.I0(shift_carry), .I1(n5), .I2(\alu_mux_sel_value[1] ), 
            .I3(alu_mux_sel_value_0__N_184), .O(n4_adj_807));   // src/flags.vhd(230[3] 234[119])
    defparam i1_4_lut_adj_273.LUT_INIT = 16'heeec;
    SB_LUT4 i2_4_lut (.I0(\instruction[14] ), .I1(n4_adj_807), .I2(arith_logical_sel_2__N_179), 
            .I3(parity), .O(carry_flag_value));   // src/flags.vhd(230[3] 234[119])
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut (.I0(flag_enable), .I1(internal_reset), .I2(wea[0]), 
            .I3(wea[0]), .O(n761));   // src/flags.vhd(91[9] 99[16])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7728_2_lut (.I0(alu_result[5]), .I1(alu_result[4]), .I2(wea[0]), 
            .I3(wea[0]), .O(n8787));
    defparam i7728_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7724_2_lut (.I0(alu_result[6]), .I1(alu_result[0]), .I2(wea[0]), 
            .I3(wea[0]), .O(n8783));
    defparam i7724_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7732_4_lut (.I0(alu_result[1]), .I1(alu_result[2]), .I2(alu_result[7]), 
            .I3(n8787), .O(n8791));
    defparam i7732_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(\instruction[15] ), .I1(\instruction[16] ), .I2(\instruction[14] ), 
            .I3(wea[0]), .O(upper_zero_sel));   // src/flags.vhd(350[20] 352[37])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i10090_4_lut (.I0(alu_result[3]), .I1(n8783), .I2(use_zero_flag), 
            .I3(zero_flag), .O(n11087));   // src/flags.vhd(357[9] 364[18])
    defparam i10090_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 carry_middle_zero_I_0_4_lut (.I0(shadow_zero_flag), .I1(n11087), 
            .I2(upper_zero_sel), .I3(n8791), .O(zero_flag_value));   // src/flags.vhd(357[9] 364[18])
    defparam carry_middle_zero_I_0_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10104_2_lut (.I0(\arith_logical_sel[0] ), .I1(\arith_logical_sel[2] ), 
            .I2(wea[0]), .I3(wea[0]), .O(n11163));   // src/zipi8.vhd(312[12:27])
    defparam i10104_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3537_4_lut (.I0(n11163), .I1(n11080), .I2(\register_vector[9] ), 
            .I3(n338), .O(n3783));   // src/zipi8.vhd(312[12:27])
    defparam i3537_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i10057_4_lut (.I0(n4), .I1(\arith_logical_sel[2] ), .I2(\register_vector[9] ), 
            .I3(\arith_logical_sel[0] ), .O(n11084));   // src/zipi8.vhd(39[28:35])
    defparam i10057_4_lut.LUT_INIT = 16'he0ac;
    SB_LUT4 i3538_3_lut (.I0(n11084), .I1(n3783), .I2(\port_id[1] ), .I3(wea[0]), 
            .O(\half_arith_logical[1] ));   // src/zipi8.vhd(39[28:35])
    defparam i3538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20_3_lut (.I0(\instruction[13] ), .I1(\instruction[14] ), .I2(\instruction[15] ), 
            .I3(wea[0]), .O(n7));
    defparam i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(carry_flag_value_N_436), .I1(\instruction[16] ), 
            .I2(n7), .I3(wea[0]), .O(\arith_logical_sel[0] ));
    defparam i1_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i602_3_lut (.I0(\instruction[16] ), .I1(\instruction[15] ), 
            .I2(\instruction[14] ), .I3(wea[0]), .O(n207));   // src/flags.vhd(302[3] 303[103])
    defparam i602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_274 (.I0(\instruction[16] ), .I1(\sx[7] ), .I2(\register_vector[8] ), 
            .I3(\instruction[3] ), .O(n687));   // src/flags.vhd(193[4:59])
    defparam i1_4_lut_adj_274.LUT_INIT = 16'ha088;
    SB_LUT4 i450_3_lut (.I0(shadow_carry_flag), .I1(\instruction[7] ), .I2(\instruction[16] ), 
            .I3(wea[0]), .O(shift_carry_value_N_413));   // src/flags.vhd(190[3] 191[51])
    defparam i450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 port_id_5__bdd_4_lut_11768 (.I0(\port_id[5] ), .I1(n722), .I2(n11107), 
            .I3(\sx[5] ), .O(n12779));
    defparam port_id_5__bdd_4_lut_11768.LUT_INIT = 16'he4aa;
    SB_LUT4 n12779_bdd_4_lut (.I0(n12779), .I1(n11109), .I2(n350), .I3(\sx[5] ), 
            .O(\half_arith_logical[5] ));
    defparam n12779_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i601_3_lut_4_lut (.I0(\instruction[16] ), .I1(\instruction[15] ), 
            .I2(carry_flag_value_N_436), .I3(arith_carry), .O(n5));   // src/flags.vhd(230[3] 234[119])
    defparam i601_3_lut_4_lut.LUT_INIT = 16'hf088;
    SB_LUT4 i2_4_lut_4_lut (.I0(arith_logical_result[7]), .I1(arith_logical_result[6]), 
            .I2(arith_logical_result[4]), .I3(arith_logical_result[5]), 
            .O(n8718));   // src/flags.vhd(147[9] 178[178])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h9661;
    SB_LUT4 i2_2_lut_4_lut (.I0(arith_logical_result[5]), .I1(arith_logical_result[7]), 
            .I2(arith_logical_result[6]), .I3(arith_logical_result[4]), 
            .O(n8728));   // src/flags.vhd(147[9] 178[178])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6986;
    SB_LUT4 i1_4_lut_4_lut (.I0(arith_logical_result[7]), .I1(arith_logical_result[6]), 
            .I2(arith_logical_result[4]), .I3(n55), .O(n4_c));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0804;
    SB_LUT4 i1_4_lut_adj_275 (.I0(\arith_logical_sel[2] ), .I1(\arith_logical_sel[0] ), 
            .I2(\sx[5] ), .I3(n338), .O(n4_adj_2));   // src/flags.vhd(67[12:28])
    defparam i1_4_lut_adj_275.LUT_INIT = 16'h3f31;
    
endmodule
//
// Verilog Description of module decode4alu
//

module decode4alu (alu_mux_sel_value, alu_mux_sel, CLK_3P3_MHZ_c, \instruction[16] , 
            \instruction[15] , \instruction[14] , carry_flag_value_N_436, 
            wea, alu_mux_sel_value_0__N_184, arith_logical_sel, n350, 
            n4247, arith_logical_sel_2__N_179, n722, \instruction[13] , 
            \sx[5] , n338, n11109);
    output [1:0]alu_mux_sel_value;
    output [1:0]alu_mux_sel;
    input CLK_3P3_MHZ_c;
    input \instruction[16] ;
    input \instruction[15] ;
    input \instruction[14] ;
    output carry_flag_value_N_436;
    input [0:0]wea;
    output alu_mux_sel_value_0__N_184;
    output [2:0]arith_logical_sel;
    output n350;
    input n4247;
    output arith_logical_sel_2__N_179;
    output n722;
    input \instruction[13] ;
    input \sx[5] ;
    input n338;
    output n11109;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [1:0]alu_mux_sel_value_c;   // src/decode4alu.vhd(48[12:29])
    
    SB_DFF alu_mux_sel_i1 (.Q(alu_mux_sel[1]), .C(CLK_3P3_MHZ_c), .D(alu_mux_sel_value[1]));   // src/decode4alu.vhd(53[9] 55[16])
    SB_LUT4 carry_flag_value_I_207_2_lut_3_lut (.I0(\instruction[16] ), .I1(\instruction[15] ), 
            .I2(\instruction[14] ), .I3(wea[0]), .O(carry_flag_value_N_436));   // src/decode4alu.vhd(71[38] 72[66])
    defparam carry_flag_value_I_207_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 alu_mux_sel_value_0__I_64_2_lut_3_lut (.I0(\instruction[16] ), 
            .I1(\instruction[15] ), .I2(\instruction[14] ), .I3(wea[0]), 
            .O(alu_mux_sel_value_0__N_184));   // src/decode4alu.vhd(71[38] 72[66])
    defparam alu_mux_sel_value_0__I_64_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF alu_mux_sel_i0 (.Q(alu_mux_sel[0]), .C(CLK_3P3_MHZ_c), .D(alu_mux_sel_value_c[0]));   // src/decode4alu.vhd(53[9] 55[16])
    SB_LUT4 i1_2_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(wea[0]), .I3(wea[0]), .O(n350));   // src/decode4alu.vhd(139[34] 140[97])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 arith_logical_sel_2__N_173_I_0_2_lut (.I0(n4247), .I1(\instruction[14] ), 
            .I2(wea[0]), .I3(wea[0]), .O(arith_logical_sel[1]));   // src/decode4alu.vhd(127[34:136])
    defparam arith_logical_sel_2__N_173_I_0_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i127_3_lut (.I0(\instruction[16] ), .I1(\instruction[14] ), 
            .I2(\instruction[15] ), .I3(wea[0]), .O(arith_logical_sel[2]));   // src/decode4alu.vhd(139[34] 140[97])
    defparam i127_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 instruction_16_downto_13_16__N_175_I_0_2_lut (.I0(\instruction[16] ), 
            .I1(\instruction[15] ), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_sel_2__N_179));   // src/decode4alu.vhd(100[34:99])
    defparam instruction_16_downto_13_16__N_175_I_0_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 arith_logical_sel_2__N_179_I_0_2_lut (.I0(arith_logical_sel_2__N_179), 
            .I1(\instruction[14] ), .I2(wea[0]), .I3(wea[0]), .O(alu_mux_sel_value[1]));   // src/decode4alu.vhd(100[34:136])
    defparam arith_logical_sel_2__N_179_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7621_2_lut_3_lut_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(n4247), .I3(\instruction[14] ), .O(n722));   // src/decode4alu.vhd(139[34] 140[97])
    defparam i7621_2_lut_3_lut_3_lut_4_lut.LUT_INIT = 16'h8d88;
    SB_LUT4 i67_3_lut (.I0(alu_mux_sel_value_0__N_184), .I1(alu_mux_sel_value[1]), 
            .I2(\instruction[13] ), .I3(wea[0]), .O(alu_mux_sel_value_c[0]));   // src/decode4alu.vhd(67[33] 74[67])
    defparam i67_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10061_2_lut_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(\sx[5] ), .I3(n338), .O(n11109));   // src/decode4alu.vhd(139[34] 140[97])
    defparam i10061_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfb9;
    
endmodule
//
// Verilog Description of module decode4_strobes_enables
//

module decode4_strobes_enables (flag_enable, CLK_3P3_MHZ_c, t_state_1_N_95, 
            register_enable, spm_enable, instruction_13_N_701, \instruction[17] , 
            \instruction[15] , \instruction[14] , flag_enable_type_N_222, 
            wea, carry_flag, pc_move_is_valid_o_N_132, \t_state[1] , 
            arith_logical_sel_2__N_179, \instruction[16] , flag_enable_type_N_216, 
            n4247, n4283, \instruction[12] , \instruction[13] , flag_enable_type_N_217);
    output flag_enable;
    input CLK_3P3_MHZ_c;
    input t_state_1_N_95;
    output register_enable;
    output spm_enable;
    input instruction_13_N_701;
    input \instruction[17] ;
    input \instruction[15] ;
    input \instruction[14] ;
    output flag_enable_type_N_222;
    input [0:0]wea;
    input carry_flag;
    output pc_move_is_valid_o_N_132;
    input \t_state[1] ;
    input arith_logical_sel_2__N_179;
    input \instruction[16] ;
    output flag_enable_type_N_216;
    output n4247;
    input n4283;
    input \instruction[12] ;
    input \instruction[13] ;
    output flag_enable_type_N_217;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    wire n498, n504, spm_enable_value_N_245, n4308, n317, n866, 
        n633, n8729;
    
    SB_DFFSR flag_enable_98 (.Q(flag_enable), .C(CLK_3P3_MHZ_c), .D(n498), 
            .R(t_state_1_N_95));   // src/decode4_strobes_enables.vhd(63[9] 81[16])
    SB_DFFSR register_enable_97 (.Q(register_enable), .C(CLK_3P3_MHZ_c), 
            .D(n504), .R(t_state_1_N_95));   // src/decode4_strobes_enables.vhd(63[9] 81[16])
    SB_DFFSR spm_enable_100 (.Q(spm_enable), .C(CLK_3P3_MHZ_c), .D(spm_enable_value_N_245), 
            .R(instruction_13_N_701));   // src/decode4_strobes_enables.vhd(63[9] 81[16])
    SB_LUT4 flag_enable_type_I_80_2_lut_3_lut (.I0(\instruction[17] ), .I1(\instruction[15] ), 
            .I2(\instruction[14] ), .I3(wea[0]), .O(flag_enable_type_N_222));   // src/decode4_strobes_enables.vhd(97[8:69])
    defparam flag_enable_type_I_80_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut (.I0(\instruction[17] ), .I1(\instruction[15] ), 
            .I2(carry_flag), .I3(wea[0]), .O(pc_move_is_valid_o_N_132));   // src/decode4_strobes_enables.vhd(97[8:69])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i3_4_lut (.I0(\t_state[1] ), .I1(\instruction[14] ), .I2(arith_logical_sel_2__N_179), 
            .I3(\instruction[17] ), .O(spm_enable_value_N_245));   // src/decode4_strobes_enables.vhd(151[22:113])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 instruction_17_downto_12_16__I_0_2_lut (.I0(\instruction[16] ), 
            .I1(\instruction[15] ), .I2(wea[0]), .I3(wea[0]), .O(flag_enable_type_N_216));   // src/decode4_strobes_enables.vhd(95[8:69])
    defparam instruction_17_downto_12_16__I_0_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4008_2_lut (.I0(\instruction[16] ), .I1(\instruction[15] ), 
            .I2(wea[0]), .I3(wea[0]), .O(n4247));
    defparam i4008_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4068_3_lut (.I0(\instruction[17] ), .I1(\instruction[15] ), 
            .I2(\instruction[14] ), .I3(wea[0]), .O(n4308));
    defparam i4068_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut (.I0(n4308), .I1(n317), .I2(n4247), .I3(n4283), 
            .O(n504));   // src/decode4_strobes_enables.vhd(130[27] 131[78])
    defparam i1_4_lut.LUT_INIT = 16'h444c;
    SB_LUT4 flag_enable_value_I_84_2_lut (.I0(\instruction[17] ), .I1(\instruction[12] ), 
            .I2(wea[0]), .I3(wea[0]), .O(n317));   // src/decode4_strobes_enables.vhd(119[23] 120[73])
    defparam flag_enable_value_I_84_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i618_4_lut (.I0(\instruction[16] ), .I1(\instruction[17] ), 
            .I2(\instruction[15] ), .I3(\instruction[14] ), .O(n866));   // src/decode4_strobes_enables.vhd(92[22] 97[144])
    defparam i618_4_lut.LUT_INIT = 16'ha022;
    SB_LUT4 i1_4_lut_adj_271 (.I0(\instruction[13] ), .I1(\instruction[14] ), 
            .I2(flag_enable_type_N_222), .I3(\instruction[17] ), .O(n633));   // src/decode4_strobes_enables.vhd(97[8:143])
    defparam i1_4_lut_adj_271.LUT_INIT = 16'h5054;
    SB_LUT4 i2_4_lut (.I0(\instruction[14] ), .I1(\instruction[16] ), .I2(flag_enable_type_N_217), 
            .I3(\instruction[17] ), .O(n8729));
    defparam i2_4_lut.LUT_INIT = 16'h0032;
    SB_LUT4 i1_4_lut_adj_272 (.I0(n8729), .I1(n317), .I2(n633), .I3(n866), 
            .O(n498));   // src/decode4_strobes_enables.vhd(119[23] 120[73])
    defparam i1_4_lut_adj_272.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_2_lut (.I0(\instruction[13] ), .I1(\instruction[15] ), .I2(wea[0]), 
            .I3(wea[0]), .O(flag_enable_type_N_217));   // src/decode4_strobes_enables.vhd(96[8:147])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    
endmodule
//
// Verilog Description of module decode4_pc_statck
//

module decode4_pc_statck (\instruction[15] , pc_mode_2__N_104, \instruction[14] , 
            \instruction[12] , n6, regbank_type_N_77, \pc_mode_2__N_158[2] , 
            pop_stack_N_164, push_stack_N_165, wea, pop_stack, \instruction[17] , 
            zero_flag, pc_move_is_valid_o_N_132, flag_enable_type_N_222, 
            carry_flag, \instruction[13] , \instruction[16] , n4283, 
            \pc_mode[0] , arith_logical_sel_2__N_179);
    input \instruction[15] ;
    output pc_mode_2__N_104;
    input \instruction[14] ;
    input \instruction[12] ;
    output n6;
    input regbank_type_N_77;
    output \pc_mode_2__N_158[2] ;
    output pop_stack_N_164;
    output push_stack_N_165;
    input [0:0]wea;
    output pop_stack;
    input \instruction[17] ;
    input zero_flag;
    input pc_move_is_valid_o_N_132;
    input flag_enable_type_N_222;
    input carry_flag;
    input \instruction[13] ;
    input \instruction[16] ;
    output n4283;
    output \pc_mode[0] ;
    input arith_logical_sel_2__N_179;
    
    
    wire n4279, n4, pc_move_is_valid_o, pc_move_is_valid_o_N_120, n4_adj_805, 
        n8719, returni_type_o_N_155;
    
    SB_LUT4 pc_mode_2__I_0_3_lut_4_lut (.I0(\instruction[15] ), .I1(n4279), 
            .I2(n4), .I3(pc_move_is_valid_o), .O(pc_mode_2__N_104));
    defparam pc_mode_2__I_0_3_lut_4_lut.LUT_INIT = 16'hf100;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\instruction[15] ), .I1(n4279), .I2(\instruction[14] ), 
            .I3(\instruction[12] ), .O(n6));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_4_lut (.I0(\instruction[15] ), .I1(\instruction[12] ), 
            .I2(\instruction[14] ), .I3(regbank_type_N_77), .O(\pc_mode_2__N_158[2] ));   // src/decode4_pc_statck.vhd(140[24] 141[94])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 push_stack_I_0_2_lut (.I0(pop_stack_N_164), .I1(\instruction[12] ), 
            .I2(wea[0]), .I3(wea[0]), .O(push_stack_N_165));   // src/decode4_pc_statck.vhd(162[23:127])
    defparam push_stack_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 pop_stack_I_0_2_lut (.I0(pop_stack_N_164), .I1(\instruction[12] ), 
            .I2(wea[0]), .I3(wea[0]), .O(pop_stack));   // src/decode4_pc_statck.vhd(151[21:146])
    defparam pop_stack_I_0_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 instruction_17_downto_12_17__I_0_106_2_lut (.I0(\instruction[17] ), 
            .I1(\instruction[15] ), .I2(wea[0]), .I3(wea[0]), .O(pc_move_is_valid_o_N_120));   // src/decode4_pc_statck.vhd(71[30:95])
    defparam instruction_17_downto_12_17__I_0_106_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut (.I0(pc_move_is_valid_o_N_120), .I1(\instruction[14] ), 
            .I2(zero_flag), .I3(pc_move_is_valid_o_N_132), .O(n4_adj_805));   // src/decode4_pc_statck.vhd(70[29] 74[143])
    defparam i1_4_lut.LUT_INIT = 16'hec28;
    SB_LUT4 i1_4_lut_adj_269 (.I0(regbank_type_N_77), .I1(flag_enable_type_N_222), 
            .I2(n4_adj_805), .I3(carry_flag), .O(pc_move_is_valid_o));   // src/decode4_pc_statck.vhd(70[29] 74[143])
    defparam i1_4_lut_adj_269.LUT_INIT = 16'hfefa;
    SB_LUT4 i4039_2_lut (.I0(\instruction[12] ), .I1(\instruction[13] ), 
            .I2(wea[0]), .I3(wea[0]), .O(n4279));
    defparam i4039_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_270 (.I0(\instruction[12] ), .I1(\instruction[16] ), 
            .I2(n4283), .I3(n4279), .O(n4));   // src/decode4_pc_statck.vhd(99[21] 103[125])
    defparam i1_4_lut_adj_270.LUT_INIT = 16'h0ace;
    SB_LUT4 i2_4_lut (.I0(\instruction[15] ), .I1(\instruction[12] ), .I2(\instruction[16] ), 
            .I3(\instruction[14] ), .O(n8719));
    defparam i2_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i3_4_lut (.I0(\instruction[12] ), .I1(pc_move_is_valid_o), .I2(returni_type_o_N_155), 
            .I3(n8719), .O(\pc_mode[0] ));
    defparam i3_4_lut.LUT_INIT = 16'hff3b;
    SB_LUT4 i4043_2_lut (.I0(\instruction[13] ), .I1(\instruction[14] ), 
            .I2(wea[0]), .I3(wea[0]), .O(n4283));
    defparam i4043_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 returni_type_o_I_55_2_lut_3_lut (.I0(arith_logical_sel_2__N_179), 
            .I1(\instruction[14] ), .I2(\instruction[13] ), .I3(wea[0]), 
            .O(returni_type_o_N_155));   // src/decode4_pc_statck.vhd(85[30] 88[63])
    defparam returni_type_o_I_55_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 pc_mode_2__N_104_I_0_2_lut_2_lut (.I0(pc_mode_2__N_104), .I1(\instruction[13] ), 
            .I2(wea[0]), .I3(wea[0]), .O(pop_stack_N_164));   // src/decode4_pc_statck.vhd(151[21:113])
    defparam pc_mode_2__N_104_I_0_2_lut_2_lut.LUT_INIT = 16'h2222;
    
endmodule
//
// Verilog Description of module arith_and_logic_operations
//

module arith_and_logic_operations (arith_logical_result, CLK_3P3_MHZ_c, 
            arith_logical_sel, \register_vector[8] , n722, n4, n11080, 
            arith_carry_in, wea, \port_id[0] , \register_vector[10] , 
            \port_id[2] , \half_arith_logical[1] , \register_vector[9] , 
            \register_vector[11] , \port_id[3] , \sx[4] , \port_id[4] , 
            \sx[6] , \port_id[6] , \half_arith_logical[5] , \sx[5] , 
            \sx[7] , carry_arith_logical_7, n350, \port_id[7] , n11084, 
            n3783, \port_id[1] , n4247, \instruction[14] , n338, n4_adj_1, 
            n11107);
    output [7:0]arith_logical_result;
    input CLK_3P3_MHZ_c;
    input [2:0]arith_logical_sel;
    input \register_vector[8] ;
    input n722;
    output n4;
    output n11080;
    input arith_carry_in;
    input [0:0]wea;
    input \port_id[0] ;
    input \register_vector[10] ;
    input \port_id[2] ;
    input \half_arith_logical[1] ;
    input \register_vector[9] ;
    input \register_vector[11] ;
    input \port_id[3] ;
    input \sx[4] ;
    input \port_id[4] ;
    input \sx[6] ;
    input \port_id[6] ;
    input \half_arith_logical[5] ;
    input \sx[5] ;
    input \sx[7] ;
    output carry_arith_logical_7;
    input n350;
    input \port_id[7] ;
    input n11084;
    input n3783;
    input \port_id[1] ;
    input n4247;
    input \instruction[14] ;
    output n338;
    input n4_adj_1;
    output n11107;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    wire [7:0]arith_logical_value;   // src/arith_and_logic_operations.vhd(50[12:31])
    
    wire n11;
    wire [7:0]half_arith_logical;   // src/arith_and_logic_operations.vhd(49[12:30])
    
    wire n8630, n8658;
    wire [7:0]carry_arith_logical;   // src/arith_and_logic_operations.vhd(51[12:31])
    
    wire n25, n13, n8664, n25_adj_798, n13_adj_799, n8654, n25_adj_800, 
        n13_adj_801, n8660, n25_adj_802, n13_adj_803, n8662, n13703, 
        n11108, n8674;
    
    SB_DFF arith_logical_result_i0 (.Q(arith_logical_result[0]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[0]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_DFF arith_logical_result_i1 (.Q(arith_logical_result[1]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[1]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_DFF arith_logical_result_i2 (.Q(arith_logical_result[2]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[2]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_DFF arith_logical_result_i3 (.Q(arith_logical_result[3]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[3]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_DFF arith_logical_result_i4 (.Q(arith_logical_result[4]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[4]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_DFF arith_logical_result_i5 (.Q(arith_logical_result[5]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[5]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_DFF arith_logical_result_i6 (.Q(arith_logical_result[6]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[6]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_DFF arith_logical_result_i7 (.Q(arith_logical_result[7]), .C(CLK_3P3_MHZ_c), 
           .D(arith_logical_value[7]));   // src/arith_and_logic_operations.vhd(56[9] 58[16])
    SB_LUT4 i24_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[1]), 
            .I2(\register_vector[8] ), .I3(n722), .O(n11));
    defparam i24_3_lut_4_lut.LUT_INIT = 16'he0ef;
    SB_LUT4 i10087_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[1]), 
            .I2(arith_logical_sel[0]), .I3(n4), .O(n11080));
    defparam i10087_3_lut_4_lut.LUT_INIT = 16'hff1f;
    SB_LUT4 half_arith_logical_7__I_0_i1_2_lut (.I0(half_arith_logical[0]), 
            .I1(arith_carry_in), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_value[0]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(\register_vector[8] ), .I3(wea[0]), .O(n8630));
    defparam i1_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_4_lut (.I0(\port_id[0] ), .I1(n8630), .I2(n8658), .I3(n11), 
            .O(half_arith_logical[0]));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i1_4_lut.LUT_INIT = 16'h72fa;
    SB_LUT4 arith_carry_in_I_0_4_lut (.I0(arith_logical_sel[2]), .I1(arith_carry_in), 
            .I2(half_arith_logical[0]), .I3(\register_vector[8] ), .O(carry_arith_logical[0]));   // src/arith_and_logic_operations.vhd(331[9] 338[18])
    defparam arith_carry_in_I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i30_3_lut (.I0(n722), .I1(arith_logical_sel[0]), .I2(\register_vector[10] ), 
            .I3(wea[0]), .O(n25));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_adj_262 (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[1]), 
            .I2(arith_logical_sel[0]), .I3(\register_vector[10] ), .O(n13));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i1_4_lut_adj_262.LUT_INIT = 16'h1505;
    SB_LUT4 i10096_4_lut (.I0(n8664), .I1(n13), .I2(\port_id[2] ), .I3(n25), 
            .O(half_arith_logical[2]));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10096_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 carry_arith_logical_0__I_0_4_lut (.I0(arith_logical_sel[2]), .I1(carry_arith_logical[0]), 
            .I2(\half_arith_logical[1] ), .I3(\register_vector[9] ), .O(carry_arith_logical[1]));   // src/arith_and_logic_operations.vhd(344[9] 351[18])
    defparam carry_arith_logical_0__I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i30_3_lut_adj_263 (.I0(n722), .I1(arith_logical_sel[0]), .I2(\register_vector[11] ), 
            .I3(wea[0]), .O(n25_adj_798));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i30_3_lut_adj_263.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_adj_264 (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[1]), 
            .I2(arith_logical_sel[0]), .I3(\register_vector[11] ), .O(n13_adj_799));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i1_4_lut_adj_264.LUT_INIT = 16'h1505;
    SB_LUT4 i10101_4_lut (.I0(n8654), .I1(n13_adj_799), .I2(\port_id[3] ), 
            .I3(n25_adj_798), .O(half_arith_logical[3]));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10101_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 carry_arith_logical_1__I_0_4_lut (.I0(arith_logical_sel[2]), .I1(carry_arith_logical[1]), 
            .I2(half_arith_logical[2]), .I3(\register_vector[10] ), .O(carry_arith_logical[2]));   // src/arith_and_logic_operations.vhd(357[9] 364[18])
    defparam carry_arith_logical_1__I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i30_3_lut_adj_265 (.I0(n722), .I1(arith_logical_sel[0]), .I2(\sx[4] ), 
            .I3(wea[0]), .O(n25_adj_800));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i30_3_lut_adj_265.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_adj_266 (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[1]), 
            .I2(arith_logical_sel[0]), .I3(\sx[4] ), .O(n13_adj_801));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i1_4_lut_adj_266.LUT_INIT = 16'h1505;
    SB_LUT4 i10099_4_lut (.I0(n8660), .I1(n13_adj_801), .I2(\port_id[4] ), 
            .I3(n25_adj_800), .O(half_arith_logical[4]));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10099_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 carry_arith_logical_2__I_0_4_lut (.I0(arith_logical_sel[2]), .I1(carry_arith_logical[2]), 
            .I2(half_arith_logical[3]), .I3(\register_vector[11] ), .O(carry_arith_logical[3]));   // src/arith_and_logic_operations.vhd(370[9] 377[18])
    defparam carry_arith_logical_2__I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 carry_arith_logical_3__I_0_4_lut (.I0(arith_logical_sel[2]), .I1(carry_arith_logical[3]), 
            .I2(half_arith_logical[4]), .I3(\sx[4] ), .O(carry_arith_logical[4]));   // src/arith_and_logic_operations.vhd(383[9] 390[18])
    defparam carry_arith_logical_3__I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i30_3_lut_adj_267 (.I0(n722), .I1(arith_logical_sel[0]), .I2(\sx[6] ), 
            .I3(wea[0]), .O(n25_adj_802));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i30_3_lut_adj_267.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_adj_268 (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[1]), 
            .I2(arith_logical_sel[0]), .I3(\sx[6] ), .O(n13_adj_803));   // src/arith_and_logic_operations.vhd(318[13] 321[94])
    defparam i1_4_lut_adj_268.LUT_INIT = 16'h1505;
    SB_LUT4 i10098_4_lut (.I0(n8662), .I1(n13_adj_803), .I2(\port_id[6] ), 
            .I3(n25_adj_802), .O(half_arith_logical[6]));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10098_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 carry_arith_logical_4__I_0_4_lut (.I0(arith_logical_sel[2]), .I1(carry_arith_logical[4]), 
            .I2(\half_arith_logical[5] ), .I3(\sx[5] ), .O(carry_arith_logical[5]));   // src/arith_and_logic_operations.vhd(396[9] 403[18])
    defparam carry_arith_logical_4__I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 carry_arith_logical_5__I_0_4_lut (.I0(arith_logical_sel[2]), .I1(carry_arith_logical[5]), 
            .I2(half_arith_logical[6]), .I3(\sx[6] ), .O(carry_arith_logical[6]));   // src/arith_and_logic_operations.vhd(409[9] 416[18])
    defparam carry_arith_logical_5__I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 carry_arith_logical_6__I_0_4_lut (.I0(arith_logical_sel[2]), .I1(carry_arith_logical[6]), 
            .I2(half_arith_logical[7]), .I3(\sx[7] ), .O(carry_arith_logical_7));   // src/arith_and_logic_operations.vhd(422[9] 429[18])
    defparam carry_arith_logical_6__I_0_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 n13703_bdd_4_lut (.I0(n13703), .I1(n11108), .I2(n350), .I3(\sx[7] ), 
            .O(half_arith_logical[7]));
    defparam n13703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 port_id_7__bdd_4_lut (.I0(\port_id[7] ), .I1(n722), .I2(n8674), 
            .I3(\sx[7] ), .O(n13703));
    defparam port_id_7__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 half_arith_logical_7__I_0_i2_2_lut_4_lut (.I0(n11084), .I1(n3783), 
            .I2(\port_id[1] ), .I3(carry_arith_logical[0]), .O(arith_logical_value[1]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(n4247), 
            .I2(\instruction[14] ), .I3(\port_id[0] ), .O(n4));   // src/arith_and_logic_operations.vhd(322[14:93])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i10095_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(n722), .I3(\sx[6] ), .O(n8662));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10095_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 and_394_i8_2_lut_3_lut (.I0(arith_logical_sel[2]), .I1(n4247), 
            .I2(\instruction[14] ), .I3(wea[0]), .O(n338));   // src/arith_and_logic_operations.vhd(321[14:63])
    defparam and_394_i8_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i10094_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(n722), .I3(\sx[4] ), .O(n8660));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10094_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 i10091_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(n722), .I3(\register_vector[11] ), .O(n8654));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10091_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 i10097_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(n722), .I3(\register_vector[10] ), .O(n8664));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10097_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 i10093_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(arith_logical_sel[0]), 
            .I2(n722), .I3(\register_vector[8] ), .O(n8658));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10093_3_lut_4_lut.LUT_INIT = 16'hf022;
    SB_LUT4 half_arith_logical_7__I_0_i3_2_lut (.I0(half_arith_logical[2]), 
            .I1(carry_arith_logical[1]), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_value[2]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 half_arith_logical_7__I_0_i4_2_lut (.I0(half_arith_logical[3]), 
            .I1(carry_arith_logical[2]), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_value[3]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 half_arith_logical_7__I_0_i5_2_lut (.I0(half_arith_logical[4]), 
            .I1(carry_arith_logical[3]), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_value[4]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 half_arith_logical_7__I_0_i6_2_lut (.I0(\half_arith_logical[5] ), 
            .I1(carry_arith_logical[4]), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_value[5]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 half_arith_logical_7__I_0_i7_2_lut (.I0(half_arith_logical[6]), 
            .I1(carry_arith_logical[5]), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_value[6]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 half_arith_logical_7__I_0_i8_2_lut (.I0(half_arith_logical[7]), 
            .I1(carry_arith_logical[6]), .I2(wea[0]), .I3(wea[0]), .O(arith_logical_value[7]));   // src/arith_and_logic_operations.vhd(441[31:79])
    defparam half_arith_logical_7__I_0_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10077_2_lut_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(n4247), 
            .I2(\instruction[14] ), .I3(n4_adj_1), .O(n11107));
    defparam i10077_2_lut_3_lut_4_lut.LUT_INIT = 16'hff45;
    SB_LUT4 i7633_2_lut_3_lut_4_lut (.I0(arith_logical_sel[2]), .I1(n4247), 
            .I2(\instruction[14] ), .I3(arith_logical_sel[0]), .O(n8674));
    defparam i7633_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ff;
    SB_LUT4 i10059_3_lut (.I0(arith_logical_sel[2]), .I1(n722), .I2(arith_logical_sel[0]), 
            .I3(wea[0]), .O(n11108));   // src/arith_and_logic_operations.vhd(318[13] 325[90])
    defparam i10059_3_lut.LUT_INIT = 16'hcdcd;
    
endmodule
//
// Verilog Description of module program_memory
//

module program_memory (wea, VCC_net, CLK_3P3_MHZ_c, bram_enable, \address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] , instruction);
    input [0:0]wea;
    input VCC_net;
    input CLK_3P3_MHZ_c;
    input bram_enable;
    input \address[10] ;
    input \address[9] ;
    input \address[8] ;
    input \address[7] ;
    input \address[6] ;
    input \address[5] ;
    input \address[4] ;
    input \address[3] ;
    input \address[2] ;
    input \address[1] ;
    input \address[0] ;
    output [17:0]instruction;
    
    wire CLK_3P3_MHZ_c /* synthesis is_clock=1 */ ;   // src/top.vhd(36[9:20])
    
    SB_RAM2048x2 Ram2048x2_inst1 (.RDATA({instruction[3:2]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst1.INIT_0 = 0000001000100100001001011111000101000101100000000000011100000010001101000111110011010110110011000000110011010100010110010100011000001011001011101110001111111111101010100101010100000000111111101010100101010100000000111010111011000000101000000000001001010101;
    defparam Ram2048x2_inst1.INIT_1 = 0001000000110000000000000011000000000000010000000000111000000001001100001000011000100110111001000000111011111111000010001000010000001110111001100010011011111111000010101010101010101000101010101000001000000000101010110000000000000000000000000000101000010011;
    defparam Ram2048x2_inst1.INIT_2 = 0101010000100000110001010101000000000101010100000000110000010101010000000000000010110001001000000000000000001100101100010010000111001100000001111001011010010000100010100110110001000100010001000100010001000100010100000101000001010000010100000001000000000100;
    defparam Ram2048x2_inst1.INIT_3 = 0000000111000101000001011010000101010100000000111111111010100001000010001111110010000000000010001100010101010000000011111111101010101011000101010100000000111111111010101011000101010100000000010101010000000000000001100100000000000010001100010101010000000001;
    defparam Ram2048x2_inst1.INIT_4 = 0011000000000000000000111111111111110000000000000000000000011111000011111100110010000100110000110011000000000100101100001111101010100101110000110010001010101010101011110000101010101010101101001000001001000000001000100000010010001111100101101000010000000000;
    defparam Ram2048x2_inst1.INIT_5 = 0000001100000000000000000000000000000000001100111000000100001100000100000001101010101000010101010000000011111111111111101010101111111010101000010101010000000000001111101010100101000000001111111110000000000001010101001100110000000000000001110001000100011100;
    defparam Ram2048x2_inst1.INIT_6 = 0101010000000011000011000001100010011000101011101110111011111111111111111101010101000000001100110000001110101010011111111110100100111000110011001001011011101110111011111000001000100010000000111111110101010100001000110000000000001010101011101110111011110010;
    defparam Ram2048x2_inst1.INIT_7 = 0101000000000000000011111111111111000100000000111111111000000000000000001111111111111100110010001000100010001000101011111111111111111111111010101111000011101000100010001000101111111111111111111111111010100011001110101000100110001001100010111111111111111101;
    defparam Ram2048x2_inst1.INIT_8 = 1111001100000011110000000000000000010010110011001010000110110010100000101100101000101011001010000010110010100010101100011000010110111101010101001100111111001111110011000000110011001111000010100000110011000000110010101010101010110011001100110000111110101010;
    defparam Ram2048x2_inst1.INIT_9 = 0000000000000000000101010100000000100000000000000000000100001100000000000001011011000000000000010000000000000101010100000000000000111110100000101000000011111111100000001111010100000101001110101010010100111111001110101011110110110000110000001110101010101010;
    defparam Ram2048x2_inst1.INIT_A = 0101010000000011111010101001000000000000001111101010100111111010101001010101000000000100000000000000000000000000000101001111101010100101010100000000111010101001010000001010101010101111001101111010101001010000111110101010010101010000000000001111111110000000;
    defparam Ram2048x2_inst1.INIT_B = 1100011000010101111101010101000000000101010100000000000000101100000000110011001110001011100100000100010000001011001100100001000010100000110000010110100000000000000100100000111010101001011010101010101111101010100101010101000000000000000000000001010100000000;
    defparam Ram2048x2_inst1.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100001100101000011011001010000010110010100010101100101000001011001010001010;
    defparam Ram2048x2_inst1.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst1.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst1.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst0 (.RDATA({instruction[1:0]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst0.INIT_0 = 0001010100000000000101001101001101100100000001010100100111001111001100000101111100011110011000111011001001000100000100000100000111000010001001001011010111000100111001001110010011100100100100111001001110010011100100001110100101100011000000110000001100000000;
    defparam Ram2048x2_inst0.INIT_1 = 0000000010110010011100001011100010010000010001000100010000000010001101010000111000011110110011100001111010101010000000000000111000011110110011100001111010101010000000000011001100100010001100110100010000000000001000010000000101000001010001110001010000110010;
    defparam Ram2048x2_inst0.INIT_2 = 1001001110000100110011100100111001001110010011100100110000111001001110010000001100111001001000000000000000000000100000100000000100001100010011000010110011111100100011100010100001001100010110000110010001110000010011000101100001100100011100000000001101000001;
    defparam Ram2048x2_inst0.INIT_3 = 0000001110011110000001001001001110010011100100111001001110001111100001000111000000000000000000001100111001001110010011100100111000010011001110010011100100111001001110010011001110010011100100111001001110000100000011001000000000000000001100111001001110010011;
    defparam Ram2048x2_inst0.INIT_4 = 1010000000000000000000111111111111110000000000000000000000111010001101101000110000111111100011011110001000111100000100000100111001001110010001010001000000000000000010000001000000000000001011000001000011000000010101110001000110001110000100100100110000000000;
    defparam Ram2048x2_inst0.INIT_5 = 0000001100000000000000000000000010010000010100010100001000001001101100000000101011111010111001001110010001110111100100111001001001001110010010111001001110010001000100111001001110001001001110010011000001101100011011001000110000000000000010110011111111111000;
    defparam Ram2048x2_inst0.INIT_6 = 1001001110010111000011010000100010001000100010001000100010111111111111111111100100111001111100110100000011100100111110010011101000110100010000001101000010001000100010110111001000010000000100111001001110010011101100110100110010001010010010001000100010110100;
    defparam Ram2048x2_inst0.INIT_7 = 1110000000000000000011111111111111001100100100111001001100000000000000001111111111111100100011011100110011001100111111111111111111111001001110011111000011010000110011001100110111111111111111111001001110010111001101001001100010001000100010011111111111111111;
    defparam Ram2048x2_inst0.INIT_8 = 1001001100000011100100000000000000100000110001000011001100010000110000000100001100010001000011001000010000110011000100001100000011110111111111001101011111001101000111000001110001010001000011100100010011000001110000000000000000100010000100100000010011100100;
    defparam Ram2048x2_inst0.INIT_9 = 0000000000000110110001101100000011000000000000000000001000011100000000000010000011000000000000100000000000001010010011100100000110100001100000011000010011100100110000101000000100000001000011100100111010100000000111101111100010100000110001001100000000000000;
    defparam Ram2048x2_inst0.INIT_A = 1001001110010001001110010011000000000000000100111001001101001110010011100100111001001001000000000000000000000000001000000100111001001110010011100100001110010011100101010000000000001011010101001110010011100000010011100100111001001110010001001110010011000000;
    defparam Ram2048x2_inst0.INIT_B = 0100001100000000110111111111000100001110010011100100000011001100000100110000000000000011010000010000000001001000001100100011110011100011110000010010010000000000001000100101001110010011100000000000001000111001001110100100111001000000000000000010010011100100;
    defparam Ram2048x2_inst0.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000001000000100001100110001000011000000010000110001000100001100100001000011001100;
    defparam Ram2048x2_inst0.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst0.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst0.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst2 (.RDATA({instruction[5:4]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst2.INIT_0 = 0000000100110000001010101000101011101000101010101010110001010000101011101010101010100100000000110001000011010001010000010000010101000000101111000011001000110101010101010101010101010101000000000000000000000000000000111111101110100010000000100000000000000000;
    defparam Ram2048x2_inst2.INIT_1 = 0100000000110100000000000011000100000000100100000000100000000000001100001111010111010100001101011101000000000000010100001111010011001100001101111111110000000000010011001101110111001111110111010100001100001000110011000001000001100000110000000000000000100011;
    defparam Ram2048x2_inst2.INIT_2 = 0000000000000000110001010101010101010000000000000000110001010101010101010000101001111110001010000000000000001101101101010000001011010010001011110010110001111101110111111011000011010100110101001101010011010100110101001101010011010100110101000000000000000000;
    defparam Ram2048x2_inst2.INIT_3 = 1110011001000000111010100101000101010101010101000000000000001011100000000111010000000001000000001100010101010101010100000000000000000011000101010101010101000000000000000011000101010101010101000000000000000010000001000100000001000000001100010101010101010100;
    defparam Ram2048x2_inst2.INIT_4 = 0010000000000000000010111111111111111000001110010011100100100110001010011000010000101001100010100110000100100100011010101010101010101010100000101011100000000000000000110000000000000000000010001110001100111000000100110000010011111010011010010111000011100100;
    defparam Ram2048x2_inst2.INIT_5 = 0000001100000000000000000000000011000011001010101000111000000100100000000010111111111110000000000000000010001000000000000000000000000000000010000000000000000000001010101010101010001010100101010101000101010101010101101000000000000000000000101100100010001000;
    defparam Ram2048x2_inst2.INIT_6 = 0000000000000111111111000001110011011100110000000000000000101111111111110000000000000000111111110000001010101010100000000000001000000000110111001110100000000000000000110010001000100000001010010101010000000000000100000000010101001101010000000000000000110001;
    defparam Ram2048x2_inst2.INIT_7 = 1010000000000000001011111111111111101000101010010101010100000000000000101111111111111110010011001100111011001101110011111111111100000000000000000011111111000000110011001100111011111111111100000000000000001111111100001100110111101101110111001111111111110000;
    defparam Ram2048x2_inst2.INIT_8 = 0000111000101110100000000000000000001011110101010010011000011000100110000111001001010001000010010100010100100100000110001001000010110100000000111100001100111000110010110000101100001100001011111101001110110000101100000000000000000000100010011000101010101010;
    defparam Ram2048x2_inst2.INIT_9 = 0000000000010101010101010111001010010011000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000101101010010010111101001010101010000001011101000101010111010101010101000101101001011111111111011000011100000111000000000000000;
    defparam Ram2048x2_inst2.INIT_A = 0000000000000000000000000000010011100100110000000000000001010101010101010101010101010000000000000000000000000000000010000101010101010101010101010101101010101010101000000000000000000010001011101010101010100000010101010101010101010101010110100101010101000000;
    defparam Ram2048x2_inst2.INIT_B = 0101001001000010110100000000100000010101010101010100001010011100001000001011011100100011010101100101011001000011010010001011000111110000111110101001010000000000000000010000101010101010100000000000000010101010101010000000000000000100111001001101010101010101;
    defparam Ram2048x2_inst2.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010010100001001100001010010011000011000100101000111001001010001000010010000;
    defparam Ram2048x2_inst2.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst2.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst2.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst3 (.RDATA({instruction[7:6]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst3.INIT_0 = 0000010000010000000001010101000101010101000000000000000101010101000101000101010101010100000101010101011011101100101100101100101001000010100011001000001100110101010101010101010101010101010101010101010101010101010101000000000000000011000000110000001000000000;
    defparam Ram2048x2_inst3.INIT_1 = 0100000000000100000011000001000100001000111000000010110010000011001100000101011100111100000101110011110000000000011000000101011100111000000101100010100000000000010001010101010001010100010101001000000100001000010001000010000001010000000000100000100000100001;
    defparam Ram2048x2_inst3.INIT_2 = 0000000000000000110000000000000000000000000000000000110000000000000000000010000000111101011000000000000000001000101000010101010110001100010001100000010000010000000000000011010011000000110000001100000011000000110000001100000011000000110000000000000000010000;
    defparam Ram2048x2_inst3.INIT_3 = 1010101010000000000000000000000000000000000000000000000000001111111000101101111000101010101000001100000000000000000000000000000000000011000000000000000000000000000000000011000000000000000000000000000000100010000010001010101010101000001100000000000000000000;
    defparam Ram2048x2_inst3.INIT_4 = 1000100000000000000000011111111111111110011111111110101010101000000111100000011000011011001001111100100110000110000011000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000010000011111111;
    defparam Ram2048x2_inst3.INIT_5 = 1000001110000000000000000010000011000011001100111101111110001100110000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000110011000000;
    defparam Ram2048x2_inst3.INIT_6 = 0000000000001001111101000010001000100001000000000000000000011111111111110000000000000000010111010000000000000000000000000000000000000000000000100000000000000000000000010000100000001000000000000000000000000000000000000000000000100000000000000000000000010000;
    defparam Ram2048x2_inst3.INIT_7 = 0000000000000000000001111111111111111000000000000000000000000000000000000111111111111111100000000000000000000000001111111111111100000000000000001101111101000000001000000001001011111111111100000000000000001001110100000000001000000010000000101111111111110000;
    defparam Ram2048x2_inst3.INIT_8 = 0010000000100000010000000000000000001001111011000001100100110000011001001100000110010011010001100100110100011001001101000110010001111100000000010100101100000010000000000000000010000010101100000000101100000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst3.INIT_9 = 0000000000000000000000000011101100000011000000000000000000000000000000000000110000000000000000000000000000000001010101010101001111101100000010000011000000000000001110111011000000100000110000000000000011101110101000001111100011010000000000000000000000000000;
    defparam Ram2048x2_inst3.INIT_A = 0101010101010101010101010101111110101010010101010101010101010101010101010101010101010100000000000000000000000000000001000101010101010101010101010101000000000000000000000000000000000000001000000000000000000000010101010101010101010101010100000000000000000000;
    defparam Ram2048x2_inst3.INIT_B = 1101000110010000111100000000010000000000000000000000100000001100001101110010001000110001111100111100110011011010001100110001110000000000110000000000000000000000000000000000000000000000000000000000000000000000000000010101010101011111101010100101010101010101;
    defparam Ram2048x2_inst3.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101100000110010011000001100100110000011001001100000110010011010001100100;
    defparam Ram2048x2_inst3.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst3.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst3.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst4 (.RDATA({instruction[9:8]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst4.INIT_0 = 1001100101001010010101010101010101010101010101010101010101010101010101010101010101010101010000010001000000000001000001000001000010110100000000010000110010010000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000000000;
    defparam Ram2048x2_inst4.INIT_1 = 0101010010100110011110001010110110011000000000100111000101000000000000010001110011000011110001000100000101010101110100000001110011000011110001000100000101010101110000010001000100010001000100010011100000011100000100010000111011100000000001000011001010110000;
    defparam Ram2048x2_inst4.INIT_2 = 0110110001101011110000011011000110110001101100011011110001000000000000000001011001110101100110010001000100010110010110011001010101100110010101011111011111010110010110011110110000110110001101100011011000110110001101100011011000110110001101100001010110100101;
    defparam Ram2048x2_inst4.INIT_3 = 1110011010001010010010110001000001101100011011000110110001100110010110110111011011011010000100011100000110110001101100011011000110101111000001101100011011000110110001101111000001101100011011000110110001101011110001000101011010000100011100000110110001101100;
    defparam Ram2048x2_inst4.INIT_4 = 1000001110010011100100111001001110010010111110010011100100101000001011100000100000101011000010111100001000001000000000001001101100011011100100101010000001101100011011100100000110110001101110010010010010010011101000000100100000000111111011000110100011100100;
    defparam Ram2048x2_inst4.INIT_5 = 0011001011110011100100111001000010000010011000101000101000001001100001000011101001100110110110110001101100001011011011000110110110110001101100000110110001101100000001101100011011000001101100011011000111100100111001011011110100010001000100010000100010000000;
    defparam Ram2048x2_inst4.INIT_6 = 0110110001101111101011101111000000110000000001000100010001110001101100011000011011000110111110111011000001101100010001101100011010101000110011000010111011101110111011111000001100111111000001101100010001101100011010101000110011000010111011101110111011111000;
    defparam Ram2048x2_inst4.INIT_7 = 1011111001001110010011100100111001001000000110110001101111100100111001001110010011100100100000000000000000000000001101101100011011011011000110111111101011101100000000000000001101101100011011011011000110111111101110110000001100000011000000110001101100011000;
    defparam Ram2048x2_inst4.INIT_8 = 1100000101000001000111100100111001000100101010001000100001100010001000011000100010000110001000100001100010001000011000100010000100011000000000001110001110101100000001000100010000000000111110110011000001000100010000011011000110111100110000001100000110110001;
    defparam Ram2048x2_inst4.INIT_9 = 1011000100010011100100111001111110110000010001000100010001000000111001001110000000001110010011100011100100111010110001101100000100010011101110111001000110110001100010000100111011101110010001101100011000010000100010010011011110110000010100000100011011000110;
    defparam Ram2048x2_inst4.INIT_A = 1100011011000100011011000110100100111001001100011011000100011011000110110001101100010110010011100100111001001110010001100001101100011011000110110001000110110001100111100001101100011001000111000110110001101011000110110001101100011011000100011011000110110001;
    defparam Ram2048x2_inst4.INIT_B = 1000100010000110011000000000001000010000000000000000010110011100110110011001100101010110010110010110011001010101100110010101010110010001000100101100010011100100111000011011000110110001100001101100011000011011000110000110110001101001001110010000011011000110;
    defparam Ram2048x2_inst4.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111001001110010001101000100010000110001000100001100010001000011000100010000110001000100001;
    defparam Ram2048x2_inst4.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst4.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst4.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst5 (.RDATA({instruction[11:10]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst5.INIT_0 = 0101010101000101010101010101010101010101010101010101010101010101010101010101010101010101010000010001000000000010000010000010000010100001000000000100010001010000000000000000000000000000000000000000000000000000000000000000000000000000100101001001010000000000;
    defparam Ram2048x2_inst5.INIT_1 = 0101010001010101010101000101010101010100001010010101001010000000001010100001010001000001010001000100000101010101010110000001010001000001010001000100000101010101010000010001000100010001000100010010100000011000000100010000010101010000000001000001000101010000;
    defparam Ram2048x2_inst5.INIT_2 = 0000000101010101110000000000010101010000000001010101110000000000000000000000000000110000000000101010101010100000000000000000000000000000000000000000000000000000000000000000000000010101000101010001010100010101000101010001010100010101000101010001010001010101;
    defparam Ram2048x2_inst5.INIT_3 = 0000000000000000000000000000000000000001010101000000000101010001001001010001001001101010101010101100000000000101010100000000010101010111000000000001010101000000000101010111000000000001010101000000000101010101011000100010101010101010101100000000000101010100;
    defparam Ram2048x2_inst5.INIT_4 = 0010100101010100000000010101010000000000010101010100000000000000000000000000000000000000000000000000000000000000001010100010101011111111000000000000101010101011111111000000101010101111111100000000000000000000000001010000000101000011110000000000000001010101;
    defparam Ram2048x2_inst5.INIT_5 = 0000000001010001010101000000100000100000000000000000000000000010001010000000000101010101011010101111111110000101000000010101011010101111111110000000000101010100001010101011111111000000000001010101001001010101000000101001011010101010101010101001000100011010;
    defparam Ram2048x2_inst5.INIT_6 = 0000000101010001010101010100000000000000001010101010101010000000000001010100000000010101000101010101000000000001010000000001010101010100000000000001010101010101010101010100000000000101000000000001010000000001010101010100000000000001010101010101010101010100;
    defparam Ram2048x2_inst5.INIT_7 = 1111111111111010101011111111101010100000000000000101010101010101000000000101010100000000000000000000000000000000000010101011111111101010111111110001010101010100000000000000000010101011111111101010111111110001010101010000000000000000000000000000000001010100;
    defparam Ram2048x2_inst5.INIT_8 = 0101101010101010011001010101000000001001101000101001100110001010011001100010100110011000101001100110001010011001100010100110011001100010101010100110011010101001101010101010101001101001111111110101010010101010101000000000010101011101110100010100101010101111;
    defparam Ram2048x2_inst5.INIT_9 = 1010111100001001010101000000111111111000000000000000000000001010010101010000011010100101010100001001010101000000000101010110000101010111111111111101000000000101010100010101111111111111010000000001010101010101000100000111010000000010101010101000000000010101;
    defparam Ram2048x2_inst5.INIT_A = 0110101010111100000000010101010101000000000110101010111100000000010101011010101011110111111110101010010101010000000001110000000001010101101010101111000000000101010111110000000001010101000111000000000101011111000000000101010110101010111100000000010101011010;
    defparam Ram2048x2_inst5.INIT_B = 0010100110011001100010101010101000000000000000000000000000001100110100000000000011111111010100010100010001000000000000010000010000000000000000000000001001010101000000011111000000000101010000000001010100000000010101000000000101010101010000000000000000010101;
    defparam Ram2048x2_inst5.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010101010000000010100010100110011000101001100110001010011001100010100110011000101001100110;
    defparam Ram2048x2_inst5.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst5.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst5.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst6 (.RDATA({instruction[13:12]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst6.INIT_0 = 1101010101100101010101010101010101010101010101010101010101010101010101010101010101010101011010011001100000000001000001000001000001010000001000000010010001011111111111111111111111111111111111111111111111111111111111111111111111110100010101000101010010101010;
    defparam Ram2048x2_inst6.INIT_1 = 0001010101110001010101010111010001010101100001110110000100010110010101010000011001101001110001100110100100000000001001010000011001101001110001100110100100000000000100010001000100010001000100011011010001010001000100010110110101010111110101100101100101010110;
    defparam Ram2048x2_inst6.INIT_2 = 1111111111011111010111111111111111111111111111111111010111111111111111110111101111011010011001000000000000001001101001100110011010011001100110100111100111101001100111110000000100110101001101010011010100110101001101010011010100110101001101010101011001010101;
    defparam Ram2048x2_inst6.INIT_3 = 1010000000111010100011111111011111111111111111111111111111011011100111011011100111101000111111110101111111111111111111111111111101111101011111111111111111111111111111111101011111111111111111111111111111001100110110011001101000111111110101111111111111111111;
    defparam Ram2048x2_inst6.INIT_4 = 1011011111111111111101111111111111111110011010101010101000000011011000001101100111100000110110000011011001111001111111001111111111111111101101110110010000000000000000101101000000000000000000010110110110100011011001111101100111111111111111111100101110101010;
    defparam Ram2048x2_inst6.INIT_5 = 0110011001110111111111111100010110010110011001101001101001011001100001011100001111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111011111111111111111011111111111111111001100110000000000000000111100000000001101;
    defparam Ram2048x2_inst6.INIT_6 = 1111111111111011011111111110110111101101110000000000000000101111111111110111111111111111101101111111011111111111111111111111111100111101100110011111110000000000000000111111011001100111011111111111111111111111111100111101100110011111110000000000000000111111;
    defparam Ram2048x2_inst6.INIT_7 = 1111111111111111110111111111111111110001111111111111111111111111111111011111111111111111000111011101110111011101111011111111111101111111111111111011011111111101110111011101111011111111111101111111111111111011011111111101111011011110110111101111111111110111;
    defparam Ram2048x2_inst6.INIT_8 = 0010111111001111100100000000000000000010010000000110001001000001100010010000011000100100000110001001000001100010010000011000100110010000000000001101101101111110110111111101111110011110011011111001100011111101111100000000000000000110011001100101111111111111;
    defparam Ram2048x2_inst6.INIT_9 = 0101010101111111111111111100111011110011000000000000000011011100000000000000100111000000000000000000000000000011111111111111010010000011111100111100111111111111111001100000111111001111001111111111111110000010011011111001000000000111111101111100000000000000;
    defparam Ram2048x2_inst6.INIT_A = 1111111111111111111111111111101010101010001111111111111111111111111111111111111111111001000000000000000000000000000010011111111111111111111111111111111111111111111001010000000000000010011001111111111111110101111111111111111111111111111111111111111111010101;
    defparam Ram2048x2_inst6.INIT_B = 0000011000100110010000000000000101111111111111111101111011110101011001100110011011101101101001101001100110011010011001100110100111110111011000111111110000000000000001100101111111111111110000000000000011111111111111111111111111111010101010101011111111111111;
    defparam Ram2048x2_inst6.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000000000000000000000011000100100000110001001000001100010010000011000100100000110001001;
    defparam Ram2048x2_inst6.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst6.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst6.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst7 (.RDATA({instruction[15:14]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst7.INIT_0 = 1010000011011110000000000000000000000000000000000000000000000000000000000000000000000000000001110011000000000000000000000000000000000000000000000001110000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000;
    defparam Ram2048x2_inst7.INIT_1 = 0111000111000111111101011100100111110101101100000011000000010100001110000000000000001011000000000000101101010101001000010000000000001011000000000000101101010101000100000000000000000000000000000000000000110101000000000101101000000110100110000010011110000101;
    defparam Ram2048x2_inst7.INIT_2 = 1010101010011010000111111111111111111010101010101010000111111111111111110000001010000001110111010101010101010111000111011100110001110111001100001110001110000111001110100000000100100000001000000010000000100000001000000010000000100000001000000111000110001100;
    defparam Ram2048x2_inst7.INIT_3 = 1111110000010110111110101010011111111111111111101010101010010000011110010000011110010000000010100001111111111111111110101010101001101000011111111111111111101010101010101000011111111111111111101010101010011001100000000011010000000010100001111111111111111110;
    defparam Ram2048x2_inst7.INIT_4 = 0011000000000000000000010101010101010100110000000000000000000011000000001100001110000000110000000011000011100011101100011011111111111111011010110000110101010101010101001010010101010101010100000010111100101000000111100000011110111111101010101000110111111111;
    defparam Ram2048x2_inst7.INIT_5 = 0000000111100100000000000000000000000000110111000011000111010000100100010100001111101011111111111111111111111010111111111111111010101010101010101010101010101001011010101010101010011010101010101010011111111111111111011001000101010101010101101000000000001100;
    defparam Ram2048x2_inst7.INIT_6 = 1010101010100111110000101000110110001101100101010101010101011111111111111110101010101010011111001010011111111111111010101010101101001000000001111011110101010101010101001011000000011110011111111111111010101010101101001000000001111011110101010101010101001011;
    defparam Ram2048x2_inst7.INIT_7 = 1111000000000000000001010101010101010001111111111111111100000000000000000101010101010101000111011001110110011101100011111111111111101010101010100111110000101001110110011101100111111111111111101010101010100111110010101101100011011000110110001111111111111110;
    defparam Ram2048x2_inst7.INIT_8 = 0100111110101010011001010101010101010000110000000000000011000000000000110000000000001100000000000011000000000000110000000000001100110001010101000000001111101000110011110000101001111000110010100011000111110000101001010101010101010000000011001101111111111111;
    defparam Ram2048x2_inst7.INIT_9 = 0000000001111111111111111101000110100100010101010101010100000001010101010101001100010101010101010101010101010110101010101010010000000011111010101000101010101010100111000000111110101010001010101010101000000001110110100011000000000111110000101001010101010101;
    defparam Ram2048x2_inst7.INIT_A = 1010101010101011111111111111000000000000001010101010101011111111111111111111111111110110010101010101010101010101010100111010101010101010101010101010111111111111110000000101010101010101110011101010101010100000111111111111111111111111111110101010101010000000;
    defparam Ram2048x2_inst7.INIT_B = 0000000000001100110001010101000001111111111111111100000110100001000111011101110011001000000111000111011100110001110111001100001110100110100000101010100101010101010101000000111111111111110101010101010110101010101010111111111111110000000000000010101010101010;
    defparam Ram2048x2_inst7.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110010101010101010100000000000000001100000000000011000000000000110000000000001100000000000011;
    defparam Ram2048x2_inst7.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst7.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst7.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 Ram2048x2_inst8 (.RDATA({instruction[17:16]}), .RCLK(CLK_3P3_MHZ_c), 
            .RCLKE(bram_enable), .RE(VCC_net), .RADDR({\address[10] , 
            \address[9] , \address[8] , \address[7] , \address[6] , 
            \address[5] , \address[4] , \address[3] , \address[2] , 
            \address[1] , \address[0] }), .WCLK(CLK_3P3_MHZ_c), .WCLKE(bram_enable), 
            .WE(wea[0]), .WADDR({\address[10] , \address[9] , \address[8] , 
            \address[7] , \address[6] , \address[5] , \address[4] , 
            \address[3] , \address[2] , \address[1] , \address[0] }), 
            .WDATA({wea, wea})) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=58, LSE_LCOL=20, LSE_RCOL=34, LSE_LLINE=87, LSE_RLINE=87 */ ;   // src/top.vhd(87[20:34])
    defparam Ram2048x2_inst8.INIT_0 = 0101000010110000101010101010101010101010101010101010101010101010101010101010101010101010101011011101111010101000101000101000101000001010101010101011001000001010101010101010101010101010101010101010101010101010101010101010101010100010000000100000001010101010;
    defparam Ram2048x2_inst8.INIT_1 = 0010001010000010101000101000000010100010110101010110100100101010110001011000011001101101001001100110110101010101000000101000011001101101001001100110110101010101001010001000100010001000100010001001011011011010100010001011010100001010101000101101110000001011;
    defparam Ram2048x2_inst8.INIT_2 = 0000000000000000001010101010101010100000000000000000001010101010101010100000000000001011001100010101010101011100101100110011001011001100110010110000110000101100110000001010101010000000100000001000000010000000100000001000000010000000100000001010001101001000;
    defparam Ram2048x2_inst8.INIT_3 = 0101011010111111010100000000101010101010101010000000000000001000110000001000110000000000000000000010101010101010101000000000000000000000101010101010101010000000000000000000101010101010101010000000000000000000000010001100000000000000000010101010101010101000;
    defparam Ram2048x2_inst8.INIT_4 = 1010000101010101010101000000000000000011000101010101010101101010001010101000110000101010100010101010001100001100001000000010101010101010110101100011000101010101010101110101010101010101010110000011010111010101011100000101110000101010000000000010111101010101;
    defparam Ram2048x2_inst8.INIT_5 = 0010001100001001010101010101000010000011001100101100101100101001110100101110101010000010101010101010101010100000101010101010100000000000000000000000000000000011100000000000000000100000000000000000101010101010101010000000000101010101010101000010101010101000;
    defparam Ram2048x2_inst8.INIT_6 = 0000000000001101010000000010100000101000000101010101010101110000000000000000000000000000110000000000101010101010100000000000001000000000100011000010100101010101010101000010001000110000101010101010100000000000001000000000100011000010100101010101010101000010;
    defparam Ram2048x2_inst8.INIT_7 = 1010010101010101010100000000000000001010101010101010101001010101010101010000000000000000101010000010100000101000001100000000000000000000000000001101010000000010100000101000001100000000000000000000000000001100000000001000001010000010100000110000000000000000;
    defparam Ram2048x2_inst8.INIT_8 = 0110101001010000110101010101010101010011000110000110011101100001100111011000011001110110000110011101100001100111011000011001110111001001010101000000110000000010100010100101000011000011000000001100100010100101000001010101010101010010001100110010101010101010;
    defparam Ram2048x2_inst8.INIT_9 = 0000000010101010101010101000000000000000010101010101010101010001010101010101110000010101010101010101010101010100000000000000101010101010100101000010000000000000001100101010101001010000100000000000000010101011001100001101101010101010100101000001010101010101;
    defparam Ram2048x2_inst8.INIT_A = 0000000000000010101010101010010101010101010000000000000010101010101010101010101010101101010101010101010101010101010111010000000000000000000000000000101010101010101001010101010101010111001101000000000000000000101010101010101010101010101000000000000000000000;
    defparam Ram2048x2_inst8.INIT_B = 1000011001110111001001010101000010101010101010101000000000000010001100110011001010000000101100101100110011001011001100110010110000001001010101000000000101010101010110100001101010101010100101010101010100000000000000101010101010100101010101010100000000000000;
    defparam Ram2048x2_inst8.INIT_C = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101010101010101010100011000011001110110000110011101100001100111011000011001110110000110011101;
    defparam Ram2048x2_inst8.INIT_D = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst8.INIT_E = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam Ram2048x2_inst8.INIT_F = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
endmodule
